

module test
(

);

  reg CLK;
  reg RST;
  wire [32-1:0] myaxi_awaddr;
  wire [8-1:0] myaxi_awlen;
  wire [3-1:0] myaxi_awsize;
  wire [2-1:0] myaxi_awburst;
  wire [1-1:0] myaxi_awlock;
  wire [4-1:0] myaxi_awcache;
  wire [3-1:0] myaxi_awprot;
  wire [4-1:0] myaxi_awqos;
  wire [2-1:0] myaxi_awuser;
  wire myaxi_awvalid;
  reg myaxi_awready;
  wire [32-1:0] myaxi_wdata;
  wire [4-1:0] myaxi_wstrb;
  wire myaxi_wlast;
  wire myaxi_wvalid;
  reg myaxi_wready;
  reg [2-1:0] myaxi_bresp;
  reg myaxi_bvalid;
  wire myaxi_bready;
  wire [32-1:0] myaxi_araddr;
  wire [8-1:0] myaxi_arlen;
  wire [3-1:0] myaxi_arsize;
  wire [2-1:0] myaxi_arburst;
  wire [1-1:0] myaxi_arlock;
  wire [4-1:0] myaxi_arcache;
  wire [3-1:0] myaxi_arprot;
  wire [4-1:0] myaxi_arqos;
  wire [2-1:0] myaxi_aruser;
  wire myaxi_arvalid;
  reg myaxi_arready;
  reg [32-1:0] myaxi_rdata;
  reg [2-1:0] myaxi_rresp;
  reg myaxi_rlast;
  reg myaxi_rvalid;
  wire myaxi_rready;
  wire [32-1:0] memory_awaddr;
  wire [8-1:0] memory_awlen;
  wire [3-1:0] memory_awsize;
  wire [2-1:0] memory_awburst;
  wire [1-1:0] memory_awlock;
  wire [4-1:0] memory_awcache;
  wire [3-1:0] memory_awprot;
  wire [4-1:0] memory_awqos;
  wire [2-1:0] memory_awuser;
  wire memory_awvalid;
  reg memory_awready;
  wire [32-1:0] memory_wdata;
  wire [4-1:0] memory_wstrb;
  wire memory_wlast;
  wire memory_wvalid;
  reg memory_wready;
  wire [2-1:0] memory_bresp;
  reg memory_bvalid;
  wire memory_bready;
  wire [32-1:0] memory_araddr;
  wire [8-1:0] memory_arlen;
  wire [3-1:0] memory_arsize;
  wire [2-1:0] memory_arburst;
  wire [1-1:0] memory_arlock;
  wire [4-1:0] memory_arcache;
  wire [3-1:0] memory_arprot;
  wire [4-1:0] memory_arqos;
  wire [2-1:0] memory_aruser;
  wire memory_arvalid;
  reg memory_arready;
  reg [32-1:0] memory_rdata;
  wire [2-1:0] memory_rresp;
  reg memory_rlast;
  reg memory_rvalid;
  wire memory_rready;
  assign memory_bresp = 0;
  assign memory_rresp = 0;
  reg [32-1:0] _memory_waddr_fsm;
  localparam _memory_waddr_fsm_init = 0;
  reg [32-1:0] _memory_wdata_fsm;
  localparam _memory_wdata_fsm_init = 0;
  reg [32-1:0] _memory_raddr_fsm;
  localparam _memory_raddr_fsm_init = 0;
  reg [32-1:0] _memory_rdata_fsm;
  localparam _memory_rdata_fsm_init = 0;
  wire _memory_wreq_fifo_enq;
  wire [41-1:0] _memory_wreq_fifo_wdata;
  wire _memory_wreq_fifo_full;
  wire _memory_wreq_fifo_almost_full;
  wire _memory_wreq_fifo_deq;
  wire [41-1:0] _memory_wreq_fifo_rdata;
  wire _memory_wreq_fifo_empty;
  wire _memory_wreq_fifo_almost_empty;

  _memory_wreq_fifo
  inst__memory_wreq_fifo
  (
    .CLK(CLK),
    .RST(RST),
    ._memory_wreq_fifo_enq(_memory_wreq_fifo_enq),
    ._memory_wreq_fifo_wdata(_memory_wreq_fifo_wdata),
    ._memory_wreq_fifo_full(_memory_wreq_fifo_full),
    ._memory_wreq_fifo_almost_full(_memory_wreq_fifo_almost_full),
    ._memory_wreq_fifo_deq(_memory_wreq_fifo_deq),
    ._memory_wreq_fifo_rdata(_memory_wreq_fifo_rdata),
    ._memory_wreq_fifo_empty(_memory_wreq_fifo_empty),
    ._memory_wreq_fifo_almost_empty(_memory_wreq_fifo_almost_empty)
  );

  reg [4-1:0] count__memory_wreq_fifo;
  wire _memory_rreq_fifo_enq;
  wire [41-1:0] _memory_rreq_fifo_wdata;
  wire _memory_rreq_fifo_full;
  wire _memory_rreq_fifo_almost_full;
  wire _memory_rreq_fifo_deq;
  wire [41-1:0] _memory_rreq_fifo_rdata;
  wire _memory_rreq_fifo_empty;
  wire _memory_rreq_fifo_almost_empty;

  _memory_rreq_fifo
  inst__memory_rreq_fifo
  (
    .CLK(CLK),
    .RST(RST),
    ._memory_rreq_fifo_enq(_memory_rreq_fifo_enq),
    ._memory_rreq_fifo_wdata(_memory_rreq_fifo_wdata),
    ._memory_rreq_fifo_full(_memory_rreq_fifo_full),
    ._memory_rreq_fifo_almost_full(_memory_rreq_fifo_almost_full),
    ._memory_rreq_fifo_deq(_memory_rreq_fifo_deq),
    ._memory_rreq_fifo_rdata(_memory_rreq_fifo_rdata),
    ._memory_rreq_fifo_empty(_memory_rreq_fifo_empty),
    ._memory_rreq_fifo_almost_empty(_memory_rreq_fifo_almost_empty)
  );

  reg [4-1:0] count__memory_rreq_fifo;
  reg [8-1:0] _memory_mem [0:2**20-1];

  initial begin
    $readmemh("memimg_parallel_add_SIMD.out", _memory_mem);
  end

  reg [33-1:0] _write_count;
  reg [32-1:0] _write_addr;
  reg [33-1:0] _read_count;
  reg [32-1:0] _read_addr;
  reg [33-1:0] _sleep_interval_count;
  reg [33-1:0] _keep_sleep_count;
  wire [32-1:0] pack_write_req_global_addr_0;
  wire [9-1:0] pack_write_req_size_1;
  assign pack_write_req_global_addr_0 = memory_awaddr;
  assign pack_write_req_size_1 = memory_awlen + 1;
  wire [41-1:0] pack_write_req_packed_2;
  assign pack_write_req_packed_2 = { pack_write_req_global_addr_0, pack_write_req_size_1 };
  assign _memory_wreq_fifo_wdata = ((_memory_waddr_fsm == 11) && memory_awvalid && memory_awready)? pack_write_req_packed_2 : 'hx;
  assign _memory_wreq_fifo_enq = ((_memory_waddr_fsm == 11) && memory_awvalid && memory_awready)? (_memory_waddr_fsm == 11) && memory_awvalid && memory_awready && !_memory_wreq_fifo_almost_full : 0;
  localparam _tmp_3 = 1;
  wire [_tmp_3-1:0] _tmp_4;
  assign _tmp_4 = !_memory_wreq_fifo_almost_full;
  reg [_tmp_3-1:0] __tmp_4_1;
  wire [32-1:0] unpack_write_req_global_addr_5;
  wire [9-1:0] unpack_write_req_size_6;
  assign unpack_write_req_global_addr_5 = _memory_wreq_fifo_rdata[40:9];
  assign unpack_write_req_size_6 = _memory_wreq_fifo_rdata[8:0];
  assign _memory_wreq_fifo_deq = ((_memory_wdata_fsm == 0) && !_memory_wreq_fifo_empty && !_memory_wreq_fifo_empty)? 1 : 0;
  wire [32-1:0] pack_read_req_global_addr_7;
  wire [9-1:0] pack_read_req_size_8;
  assign pack_read_req_global_addr_7 = memory_araddr;
  assign pack_read_req_size_8 = memory_arlen + 1;
  wire [41-1:0] pack_read_req_packed_9;
  assign pack_read_req_packed_9 = { pack_read_req_global_addr_7, pack_read_req_size_8 };
  assign _memory_rreq_fifo_wdata = ((_memory_raddr_fsm == 1) && memory_arvalid && memory_arready)? pack_read_req_packed_9 : 'hx;
  assign _memory_rreq_fifo_enq = ((_memory_raddr_fsm == 1) && memory_arvalid && memory_arready)? (_memory_raddr_fsm == 1) && memory_arvalid && memory_arready && !_memory_rreq_fifo_almost_full : 0;
  localparam _tmp_10 = 1;
  wire [_tmp_10-1:0] _tmp_11;
  assign _tmp_11 = !_memory_rreq_fifo_almost_full;
  reg [_tmp_10-1:0] __tmp_11_1;
  wire [32-1:0] unpack_read_req_global_addr_12;
  wire [9-1:0] unpack_read_req_size_13;
  assign unpack_read_req_global_addr_12 = _memory_rreq_fifo_rdata[40:9];
  assign unpack_read_req_size_13 = _memory_rreq_fifo_rdata[8:0];
  assign _memory_rreq_fifo_deq = ((_memory_rdata_fsm == 0) && !_memory_rreq_fifo_empty && !_memory_rreq_fifo_empty)? 1 : 0;
  reg [32-1:0] _d1__memory_rdata_fsm;
  reg __memory_rdata_fsm_cond_11_0_1;
  assign memory_awaddr = myaxi_awaddr;
  assign memory_awlen = myaxi_awlen;
  assign memory_awsize = myaxi_awsize;
  assign memory_awburst = myaxi_awburst;
  assign memory_awlock = myaxi_awlock;
  assign memory_awcache = myaxi_awcache;
  assign memory_awprot = myaxi_awprot;
  assign memory_awqos = myaxi_awqos;
  assign memory_awuser = myaxi_awuser;
  assign memory_awvalid = myaxi_awvalid;
  wire _tmp_14;
  assign _tmp_14 = memory_awready;

  always @(*) begin
    myaxi_awready = _tmp_14;
  end

  assign memory_wdata = myaxi_wdata;
  assign memory_wstrb = myaxi_wstrb;
  assign memory_wlast = myaxi_wlast;
  assign memory_wvalid = myaxi_wvalid;
  wire _tmp_15;
  assign _tmp_15 = memory_wready;

  always @(*) begin
    myaxi_wready = _tmp_15;
  end

  wire [2-1:0] _tmp_16;
  assign _tmp_16 = memory_bresp;

  always @(*) begin
    myaxi_bresp = _tmp_16;
  end

  wire _tmp_17;
  assign _tmp_17 = memory_bvalid;

  always @(*) begin
    myaxi_bvalid = _tmp_17;
  end

  assign memory_bready = myaxi_bready;
  assign memory_araddr = myaxi_araddr;
  assign memory_arlen = myaxi_arlen;
  assign memory_arsize = myaxi_arsize;
  assign memory_arburst = myaxi_arburst;
  assign memory_arlock = myaxi_arlock;
  assign memory_arcache = myaxi_arcache;
  assign memory_arprot = myaxi_arprot;
  assign memory_arqos = myaxi_arqos;
  assign memory_aruser = myaxi_aruser;
  assign memory_arvalid = myaxi_arvalid;
  wire _tmp_18;
  assign _tmp_18 = memory_arready;

  always @(*) begin
    myaxi_arready = _tmp_18;
  end

  wire [32-1:0] _tmp_19;
  assign _tmp_19 = memory_rdata;

  always @(*) begin
    myaxi_rdata = _tmp_19;
  end

  wire [2-1:0] _tmp_20;
  assign _tmp_20 = memory_rresp;

  always @(*) begin
    myaxi_rresp = _tmp_20;
  end

  wire _tmp_21;
  assign _tmp_21 = memory_rlast;

  always @(*) begin
    myaxi_rlast = _tmp_21;
  end

  wire _tmp_22;
  assign _tmp_22 = memory_rvalid;

  always @(*) begin
    myaxi_rvalid = _tmp_22;
  end

  assign memory_rready = myaxi_rready;

  blinkled
  uut
  (
    .CLK(CLK),
    .RST(RST),
    .myaxi_awaddr(myaxi_awaddr),
    .myaxi_awlen(myaxi_awlen),
    .myaxi_awsize(myaxi_awsize),
    .myaxi_awburst(myaxi_awburst),
    .myaxi_awlock(myaxi_awlock),
    .myaxi_awcache(myaxi_awcache),
    .myaxi_awprot(myaxi_awprot),
    .myaxi_awqos(myaxi_awqos),
    .myaxi_awuser(myaxi_awuser),
    .myaxi_awvalid(myaxi_awvalid),
    .myaxi_awready(myaxi_awready),
    .myaxi_wdata(myaxi_wdata),
    .myaxi_wstrb(myaxi_wstrb),
    .myaxi_wlast(myaxi_wlast),
    .myaxi_wvalid(myaxi_wvalid),
    .myaxi_wready(myaxi_wready),
    .myaxi_bresp(myaxi_bresp),
    .myaxi_bvalid(myaxi_bvalid),
    .myaxi_bready(myaxi_bready),
    .myaxi_araddr(myaxi_araddr),
    .myaxi_arlen(myaxi_arlen),
    .myaxi_arsize(myaxi_arsize),
    .myaxi_arburst(myaxi_arburst),
    .myaxi_arlock(myaxi_arlock),
    .myaxi_arcache(myaxi_arcache),
    .myaxi_arprot(myaxi_arprot),
    .myaxi_arqos(myaxi_arqos),
    .myaxi_aruser(myaxi_aruser),
    .myaxi_arvalid(myaxi_arvalid),
    .myaxi_arready(myaxi_arready),
    .myaxi_rdata(myaxi_rdata),
    .myaxi_rresp(myaxi_rresp),
    .myaxi_rlast(myaxi_rlast),
    .myaxi_rvalid(myaxi_rvalid),
    .myaxi_rready(myaxi_rready)
  );


  initial begin
    CLK = 0;
    forever begin
      #5 CLK = !CLK;
    end
  end


  initial begin
    RST = 0;
    memory_awready = 0;
    memory_wready = 0;
    memory_bvalid = 0;
    memory_arready = 0;
    memory_rdata = 0;
    memory_rlast = 0;
    memory_rvalid = 0;
    _memory_waddr_fsm = _memory_waddr_fsm_init;
    _memory_wdata_fsm = _memory_wdata_fsm_init;
    _memory_raddr_fsm = _memory_raddr_fsm_init;
    _memory_rdata_fsm = _memory_rdata_fsm_init;
    count__memory_wreq_fifo = 0;
    count__memory_rreq_fifo = 0;
    _write_count = 0;
    _write_addr = 0;
    _read_count = 0;
    _read_addr = 0;
    _sleep_interval_count = 0;
    _keep_sleep_count = 0;
    __tmp_4_1 = 0;
    __tmp_11_1 = 0;
    _d1__memory_rdata_fsm = _memory_rdata_fsm_init;
    __memory_rdata_fsm_cond_11_0_1 = 0;
    #100;
    RST = 1;
    #100;
    RST = 0;
    #1000000;
    $finish;
  end


  always @(posedge CLK) begin
    if(RST) begin
      _keep_sleep_count <= 0;
      _sleep_interval_count <= 0;
    end else begin
      if(_sleep_interval_count == 15) begin
        _keep_sleep_count <= _keep_sleep_count + 1;
      end 
      if((_sleep_interval_count == 15) && (_keep_sleep_count == 3)) begin
        _keep_sleep_count <= 0;
      end 
      if(_sleep_interval_count < 15) begin
        _sleep_interval_count <= _sleep_interval_count + 1;
      end 
      if((_keep_sleep_count == 3) && (_sleep_interval_count == 15)) begin
        _sleep_interval_count <= 0;
      end 
      if((_memory_wdata_fsm == 1) && memory_wvalid && memory_wready && memory_wstrb[0]) begin
        _memory_mem[_write_addr + 0] <= memory_wdata[7:0];
      end 
      if((_memory_wdata_fsm == 1) && memory_wvalid && memory_wready && memory_wstrb[1]) begin
        _memory_mem[_write_addr + 1] <= memory_wdata[15:8];
      end 
      if((_memory_wdata_fsm == 1) && memory_wvalid && memory_wready && memory_wstrb[2]) begin
        _memory_mem[_write_addr + 2] <= memory_wdata[23:16];
      end 
      if((_memory_wdata_fsm == 1) && memory_wvalid && memory_wready && memory_wstrb[3]) begin
        _memory_mem[_write_addr + 3] <= memory_wdata[31:24];
      end 
    end
  end

  localparam _memory_waddr_fsm_1 = 1;
  localparam _memory_waddr_fsm_2 = 2;
  localparam _memory_waddr_fsm_3 = 3;
  localparam _memory_waddr_fsm_4 = 4;
  localparam _memory_waddr_fsm_5 = 5;
  localparam _memory_waddr_fsm_6 = 6;
  localparam _memory_waddr_fsm_7 = 7;
  localparam _memory_waddr_fsm_8 = 8;
  localparam _memory_waddr_fsm_9 = 9;
  localparam _memory_waddr_fsm_10 = 10;
  localparam _memory_waddr_fsm_11 = 11;

  always @(posedge CLK) begin
    if(RST) begin
      _memory_waddr_fsm <= _memory_waddr_fsm_init;
      memory_awready <= 0;
    end else begin
      case(_memory_waddr_fsm)
        _memory_waddr_fsm_init: begin
          memory_awready <= 0;
          if(memory_awvalid) begin
            _memory_waddr_fsm <= _memory_waddr_fsm_1;
          end 
        end
        _memory_waddr_fsm_1: begin
          _memory_waddr_fsm <= _memory_waddr_fsm_2;
        end
        _memory_waddr_fsm_2: begin
          _memory_waddr_fsm <= _memory_waddr_fsm_3;
        end
        _memory_waddr_fsm_3: begin
          _memory_waddr_fsm <= _memory_waddr_fsm_4;
        end
        _memory_waddr_fsm_4: begin
          _memory_waddr_fsm <= _memory_waddr_fsm_5;
        end
        _memory_waddr_fsm_5: begin
          _memory_waddr_fsm <= _memory_waddr_fsm_6;
        end
        _memory_waddr_fsm_6: begin
          _memory_waddr_fsm <= _memory_waddr_fsm_7;
        end
        _memory_waddr_fsm_7: begin
          _memory_waddr_fsm <= _memory_waddr_fsm_8;
        end
        _memory_waddr_fsm_8: begin
          _memory_waddr_fsm <= _memory_waddr_fsm_9;
        end
        _memory_waddr_fsm_9: begin
          _memory_waddr_fsm <= _memory_waddr_fsm_10;
        end
        _memory_waddr_fsm_10: begin
          _memory_waddr_fsm <= _memory_waddr_fsm_11;
        end
        _memory_waddr_fsm_11: begin
          if(!_memory_wreq_fifo_almost_full) begin
            memory_awready <= 1;
          end 
          if(memory_awvalid && memory_awready) begin
            memory_awready <= 0;
          end 
          if(!memory_awvalid) begin
            _memory_waddr_fsm <= _memory_waddr_fsm_init;
          end 
          if(memory_awvalid && memory_awready) begin
            _memory_waddr_fsm <= _memory_waddr_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam _memory_wdata_fsm_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      _memory_wdata_fsm <= _memory_wdata_fsm_init;
      memory_bvalid <= 0;
      _write_addr <= 0;
      _write_count <= 0;
      memory_wready <= 0;
    end else begin
      case(_memory_wdata_fsm)
        _memory_wdata_fsm_init: begin
          memory_bvalid <= 0;
          if(!_memory_wreq_fifo_empty) begin
            _write_addr <= unpack_write_req_global_addr_5;
            _write_count <= unpack_write_req_size_6;
            memory_wready <= 1;
          end 
          if(!_memory_wreq_fifo_empty) begin
            _memory_wdata_fsm <= _memory_wdata_fsm_1;
          end 
        end
        _memory_wdata_fsm_1: begin
          if(memory_wvalid && memory_wready) begin
            _write_addr <= _write_addr + 4;
            _write_count <= _write_count - 1;
          end 
          if(_sleep_interval_count == 15) begin
            memory_wready <= 0;
          end else begin
            memory_wready <= 1;
          end
          if(memory_wvalid && memory_wready && (_write_count == 1)) begin
            memory_wready <= 0;
            memory_bvalid <= 1;
          end 
          if(memory_wvalid && memory_wready && memory_wlast) begin
            memory_wready <= 0;
            memory_bvalid <= 1;
          end 
          if(memory_wvalid && memory_wready && (_write_count == 1)) begin
            _memory_wdata_fsm <= _memory_wdata_fsm_init;
          end 
          if(memory_wvalid && memory_wready && memory_wlast) begin
            _memory_wdata_fsm <= _memory_wdata_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam _memory_raddr_fsm_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      _memory_raddr_fsm <= _memory_raddr_fsm_init;
      memory_arready <= 0;
    end else begin
      case(_memory_raddr_fsm)
        _memory_raddr_fsm_init: begin
          memory_arready <= 0;
          if(memory_arvalid) begin
            _memory_raddr_fsm <= _memory_raddr_fsm_1;
          end 
        end
        _memory_raddr_fsm_1: begin
          if(!_memory_rreq_fifo_almost_full) begin
            memory_arready <= 1;
          end 
          if(memory_arvalid && memory_arready) begin
            memory_arready <= 0;
          end 
          if(!memory_arvalid) begin
            _memory_raddr_fsm <= _memory_raddr_fsm_init;
          end 
          if(memory_arvalid && memory_arready) begin
            _memory_raddr_fsm <= _memory_raddr_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam _memory_rdata_fsm_1 = 1;
  localparam _memory_rdata_fsm_2 = 2;
  localparam _memory_rdata_fsm_3 = 3;
  localparam _memory_rdata_fsm_4 = 4;
  localparam _memory_rdata_fsm_5 = 5;
  localparam _memory_rdata_fsm_6 = 6;
  localparam _memory_rdata_fsm_7 = 7;
  localparam _memory_rdata_fsm_8 = 8;
  localparam _memory_rdata_fsm_9 = 9;
  localparam _memory_rdata_fsm_10 = 10;
  localparam _memory_rdata_fsm_11 = 11;

  always @(posedge CLK) begin
    if(RST) begin
      _memory_rdata_fsm <= _memory_rdata_fsm_init;
      _d1__memory_rdata_fsm <= _memory_rdata_fsm_init;
      _read_addr <= 0;
      _read_count <= 0;
      memory_rdata[7:0] <= (0 >> 0) & { 8{ 1'd1 } };
      memory_rdata[15:8] <= (0 >> 8) & { 8{ 1'd1 } };
      memory_rdata[23:16] <= (0 >> 16) & { 8{ 1'd1 } };
      memory_rdata[31:24] <= (0 >> 24) & { 8{ 1'd1 } };
      memory_rvalid <= 0;
      memory_rlast <= 0;
      __memory_rdata_fsm_cond_11_0_1 <= 0;
      memory_rdata <= 0;
    end else begin
      _d1__memory_rdata_fsm <= _memory_rdata_fsm;
      case(_d1__memory_rdata_fsm)
        _memory_rdata_fsm_11: begin
          if(__memory_rdata_fsm_cond_11_0_1) begin
            memory_rvalid <= 0;
            memory_rlast <= 0;
          end 
        end
      endcase
      case(_memory_rdata_fsm)
        _memory_rdata_fsm_init: begin
          if(!_memory_rreq_fifo_empty) begin
            _read_addr <= unpack_read_req_global_addr_12;
            _read_count <= unpack_read_req_size_13;
          end 
          if(!_memory_rreq_fifo_empty) begin
            _memory_rdata_fsm <= _memory_rdata_fsm_1;
          end 
        end
        _memory_rdata_fsm_1: begin
          _memory_rdata_fsm <= _memory_rdata_fsm_2;
        end
        _memory_rdata_fsm_2: begin
          _memory_rdata_fsm <= _memory_rdata_fsm_3;
        end
        _memory_rdata_fsm_3: begin
          _memory_rdata_fsm <= _memory_rdata_fsm_4;
        end
        _memory_rdata_fsm_4: begin
          _memory_rdata_fsm <= _memory_rdata_fsm_5;
        end
        _memory_rdata_fsm_5: begin
          _memory_rdata_fsm <= _memory_rdata_fsm_6;
        end
        _memory_rdata_fsm_6: begin
          _memory_rdata_fsm <= _memory_rdata_fsm_7;
        end
        _memory_rdata_fsm_7: begin
          _memory_rdata_fsm <= _memory_rdata_fsm_8;
        end
        _memory_rdata_fsm_8: begin
          _memory_rdata_fsm <= _memory_rdata_fsm_9;
        end
        _memory_rdata_fsm_9: begin
          _memory_rdata_fsm <= _memory_rdata_fsm_10;
        end
        _memory_rdata_fsm_10: begin
          _memory_rdata_fsm <= _memory_rdata_fsm_11;
        end
        _memory_rdata_fsm_11: begin
          if(memory_rready | !memory_rvalid) begin
            memory_rdata[7:0] <= _memory_mem[_read_addr + 0];
          end 
          if(memory_rready | !memory_rvalid) begin
            memory_rdata[15:8] <= _memory_mem[_read_addr + 1];
          end 
          if(memory_rready | !memory_rvalid) begin
            memory_rdata[23:16] <= _memory_mem[_read_addr + 2];
          end 
          if(memory_rready | !memory_rvalid) begin
            memory_rdata[31:24] <= _memory_mem[_read_addr + 3];
          end 
          if((_sleep_interval_count < 15) && (_read_count > 0) && memory_rready | !memory_rvalid) begin
            memory_rvalid <= 1;
            _read_addr <= _read_addr + 4;
            _read_count <= _read_count - 1;
          end 
          if((_sleep_interval_count < 15) && (_read_count == 1) && memory_rready | !memory_rvalid) begin
            memory_rlast <= 1;
          end 
          __memory_rdata_fsm_cond_11_0_1 <= 1;
          if(memory_rvalid && !memory_rready) begin
            memory_rvalid <= memory_rvalid;
            memory_rdata <= memory_rdata;
            memory_rlast <= memory_rlast;
          end 
          if(memory_rvalid && memory_rready && (_read_count == 0)) begin
            _memory_rdata_fsm <= _memory_rdata_fsm_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      count__memory_wreq_fifo <= 0;
      __tmp_4_1 <= 0;
    end else begin
      if(_memory_wreq_fifo_enq && !_memory_wreq_fifo_full && (_memory_wreq_fifo_deq && !_memory_wreq_fifo_empty)) begin
        count__memory_wreq_fifo <= count__memory_wreq_fifo;
      end else if(_memory_wreq_fifo_enq && !_memory_wreq_fifo_full) begin
        count__memory_wreq_fifo <= count__memory_wreq_fifo + 1;
      end else if(_memory_wreq_fifo_deq && !_memory_wreq_fifo_empty) begin
        count__memory_wreq_fifo <= count__memory_wreq_fifo - 1;
      end 
      __tmp_4_1 <= _tmp_4;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      count__memory_rreq_fifo <= 0;
      __tmp_11_1 <= 0;
    end else begin
      if(_memory_rreq_fifo_enq && !_memory_rreq_fifo_full && (_memory_rreq_fifo_deq && !_memory_rreq_fifo_empty)) begin
        count__memory_rreq_fifo <= count__memory_rreq_fifo;
      end else if(_memory_rreq_fifo_enq && !_memory_rreq_fifo_full) begin
        count__memory_rreq_fifo <= count__memory_rreq_fifo + 1;
      end else if(_memory_rreq_fifo_deq && !_memory_rreq_fifo_empty) begin
        count__memory_rreq_fifo <= count__memory_rreq_fifo - 1;
      end 
      __tmp_11_1 <= _tmp_11;
    end
  end


endmodule



module _memory_wreq_fifo
(
  input CLK,
  input RST,
  input _memory_wreq_fifo_enq,
  input [41-1:0] _memory_wreq_fifo_wdata,
  output _memory_wreq_fifo_full,
  output _memory_wreq_fifo_almost_full,
  input _memory_wreq_fifo_deq,
  output [41-1:0] _memory_wreq_fifo_rdata,
  output _memory_wreq_fifo_empty,
  output _memory_wreq_fifo_almost_empty
);

  reg [41-1:0] mem [0:8-1];
  reg [3-1:0] head;
  reg [3-1:0] tail;
  wire is_empty;
  wire is_almost_empty;
  wire is_full;
  wire is_almost_full;
  assign is_empty = head == tail;
  assign is_almost_empty = head == (tail + 1 & 7);
  assign is_full = (head + 1 & 7) == tail;
  assign is_almost_full = (head + 2 & 7) == tail;
  wire [41-1:0] rdata;
  assign _memory_wreq_fifo_full = is_full;
  assign _memory_wreq_fifo_almost_full = is_almost_full || is_full;
  assign _memory_wreq_fifo_empty = is_empty;
  assign _memory_wreq_fifo_almost_empty = is_almost_empty || is_empty;
  assign rdata = mem[tail];
  assign _memory_wreq_fifo_rdata = rdata;

  always @(posedge CLK) begin
    if(RST) begin
      head <= 0;
      tail <= 0;
    end else begin
      if(_memory_wreq_fifo_enq && !is_full) begin
        mem[head] <= _memory_wreq_fifo_wdata;
        head <= head + 1;
      end 
      if(_memory_wreq_fifo_deq && !is_empty) begin
        tail <= tail + 1;
      end 
    end
  end


endmodule



module _memory_rreq_fifo
(
  input CLK,
  input RST,
  input _memory_rreq_fifo_enq,
  input [41-1:0] _memory_rreq_fifo_wdata,
  output _memory_rreq_fifo_full,
  output _memory_rreq_fifo_almost_full,
  input _memory_rreq_fifo_deq,
  output [41-1:0] _memory_rreq_fifo_rdata,
  output _memory_rreq_fifo_empty,
  output _memory_rreq_fifo_almost_empty
);

  reg [41-1:0] mem [0:8-1];
  reg [3-1:0] head;
  reg [3-1:0] tail;
  wire is_empty;
  wire is_almost_empty;
  wire is_full;
  wire is_almost_full;
  assign is_empty = head == tail;
  assign is_almost_empty = head == (tail + 1 & 7);
  assign is_full = (head + 1 & 7) == tail;
  assign is_almost_full = (head + 2 & 7) == tail;
  wire [41-1:0] rdata;
  assign _memory_rreq_fifo_full = is_full;
  assign _memory_rreq_fifo_almost_full = is_almost_full || is_full;
  assign _memory_rreq_fifo_empty = is_empty;
  assign _memory_rreq_fifo_almost_empty = is_almost_empty || is_empty;
  assign rdata = mem[tail];
  assign _memory_rreq_fifo_rdata = rdata;

  always @(posedge CLK) begin
    if(RST) begin
      head <= 0;
      tail <= 0;
    end else begin
      if(_memory_rreq_fifo_enq && !is_full) begin
        mem[head] <= _memory_rreq_fifo_wdata;
        head <= head + 1;
      end 
      if(_memory_rreq_fifo_deq && !is_empty) begin
        tail <= tail + 1;
      end 
    end
  end


endmodule



module blinkled
(
  input CLK,
  input RST,
  output reg [32-1:0] myaxi_awaddr,
  output reg [8-1:0] myaxi_awlen,
  output [3-1:0] myaxi_awsize,
  output [2-1:0] myaxi_awburst,
  output [1-1:0] myaxi_awlock,
  output [4-1:0] myaxi_awcache,
  output [3-1:0] myaxi_awprot,
  output [4-1:0] myaxi_awqos,
  output [2-1:0] myaxi_awuser,
  output reg myaxi_awvalid,
  input myaxi_awready,
  output reg [32-1:0] myaxi_wdata,
  output reg [4-1:0] myaxi_wstrb,
  output reg myaxi_wlast,
  output reg myaxi_wvalid,
  input myaxi_wready,
  input [2-1:0] myaxi_bresp,
  input myaxi_bvalid,
  output myaxi_bready,
  output reg [32-1:0] myaxi_araddr,
  output reg [8-1:0] myaxi_arlen,
  output [3-1:0] myaxi_arsize,
  output [2-1:0] myaxi_arburst,
  output [1-1:0] myaxi_arlock,
  output [4-1:0] myaxi_arcache,
  output [3-1:0] myaxi_arprot,
  output [4-1:0] myaxi_arqos,
  output [2-1:0] myaxi_aruser,
  output reg myaxi_arvalid,
  input myaxi_arready,
  input [32-1:0] myaxi_rdata,
  input [2-1:0] myaxi_rresp,
  input myaxi_rlast,
  input myaxi_rvalid,
  output myaxi_rready
);

  assign myaxi_awsize = 2;
  assign myaxi_awburst = 1;
  assign myaxi_awlock = 0;
  assign myaxi_awcache = 3;
  assign myaxi_awprot = 0;
  assign myaxi_awqos = 0;
  assign myaxi_awuser = 0;
  assign myaxi_bready = 1;
  assign myaxi_arsize = 2;
  assign myaxi_arburst = 1;
  assign myaxi_arlock = 0;
  assign myaxi_arcache = 3;
  assign myaxi_arprot = 0;
  assign myaxi_arqos = 0;
  assign myaxi_aruser = 0;
  reg [3-1:0] outstanding_wcount_0;
  reg _myaxi_read_start;
  reg [8-1:0] _myaxi_read_op_sel;
  reg [32-1:0] _myaxi_read_global_addr;
  reg [33-1:0] _myaxi_read_global_size;
  reg [32-1:0] _myaxi_read_local_addr;
  reg [32-1:0] _myaxi_read_local_stride;
  reg [33-1:0] _myaxi_read_local_size;
  reg [32-1:0] _myaxi_read_local_blocksize;
  wire _myaxi_read_req_fifo_enq;
  wire [137-1:0] _myaxi_read_req_fifo_wdata;
  wire _myaxi_read_req_fifo_full;
  wire _myaxi_read_req_fifo_almost_full;
  wire _myaxi_read_req_fifo_deq;
  wire [137-1:0] _myaxi_read_req_fifo_rdata;
  wire _myaxi_read_req_fifo_empty;
  wire _myaxi_read_req_fifo_almost_empty;

  _myaxi_read_req_fifo
  inst__myaxi_read_req_fifo
  (
    .CLK(CLK),
    .RST(RST),
    ._myaxi_read_req_fifo_enq(_myaxi_read_req_fifo_enq),
    ._myaxi_read_req_fifo_wdata(_myaxi_read_req_fifo_wdata),
    ._myaxi_read_req_fifo_full(_myaxi_read_req_fifo_full),
    ._myaxi_read_req_fifo_almost_full(_myaxi_read_req_fifo_almost_full),
    ._myaxi_read_req_fifo_deq(_myaxi_read_req_fifo_deq),
    ._myaxi_read_req_fifo_rdata(_myaxi_read_req_fifo_rdata),
    ._myaxi_read_req_fifo_empty(_myaxi_read_req_fifo_empty),
    ._myaxi_read_req_fifo_almost_empty(_myaxi_read_req_fifo_almost_empty)
  );

  reg [4-1:0] count__myaxi_read_req_fifo;
  wire [8-1:0] _myaxi_read_op_sel_fifo;
  wire [32-1:0] _myaxi_read_local_addr_fifo;
  wire [32-1:0] _myaxi_read_local_stride_fifo;
  wire [33-1:0] _myaxi_read_local_size_fifo;
  wire [32-1:0] _myaxi_read_local_blocksize_fifo;
  wire [8-1:0] unpack_read_req_op_sel_1;
  wire [32-1:0] unpack_read_req_local_addr_2;
  wire [32-1:0] unpack_read_req_local_stride_3;
  wire [33-1:0] unpack_read_req_local_size_4;
  wire [32-1:0] unpack_read_req_local_blocksize_5;
  assign unpack_read_req_op_sel_1 = _myaxi_read_req_fifo_rdata[136:129];
  assign unpack_read_req_local_addr_2 = _myaxi_read_req_fifo_rdata[128:97];
  assign unpack_read_req_local_stride_3 = _myaxi_read_req_fifo_rdata[96:65];
  assign unpack_read_req_local_size_4 = _myaxi_read_req_fifo_rdata[64:32];
  assign unpack_read_req_local_blocksize_5 = _myaxi_read_req_fifo_rdata[31:0];
  assign _myaxi_read_op_sel_fifo = unpack_read_req_op_sel_1;
  assign _myaxi_read_local_addr_fifo = unpack_read_req_local_addr_2;
  assign _myaxi_read_local_stride_fifo = unpack_read_req_local_stride_3;
  assign _myaxi_read_local_size_fifo = unpack_read_req_local_size_4;
  assign _myaxi_read_local_blocksize_fifo = unpack_read_req_local_blocksize_5;
  reg [8-1:0] _myaxi_read_op_sel_buf;
  reg [32-1:0] _myaxi_read_local_addr_buf;
  reg [32-1:0] _myaxi_read_local_stride_buf;
  reg [33-1:0] _myaxi_read_local_size_buf;
  reg [32-1:0] _myaxi_read_local_blocksize_buf;
  reg _myaxi_read_req_idle;
  reg _myaxi_read_data_idle;
  wire _myaxi_read_idle;
  assign _myaxi_read_idle = !_myaxi_read_start && _myaxi_read_req_idle && _myaxi_read_req_fifo_empty && _myaxi_read_data_idle;
  reg _myaxi_write_start;
  reg [8-1:0] _myaxi_write_op_sel;
  reg [32-1:0] _myaxi_write_global_addr;
  reg [33-1:0] _myaxi_write_global_size;
  reg [32-1:0] _myaxi_write_local_addr;
  reg [32-1:0] _myaxi_write_local_stride;
  reg [33-1:0] _myaxi_write_local_size;
  reg [32-1:0] _myaxi_write_local_blocksize;
  wire _myaxi_write_req_fifo_enq;
  wire [137-1:0] _myaxi_write_req_fifo_wdata;
  wire _myaxi_write_req_fifo_full;
  wire _myaxi_write_req_fifo_almost_full;
  wire _myaxi_write_req_fifo_deq;
  wire [137-1:0] _myaxi_write_req_fifo_rdata;
  wire _myaxi_write_req_fifo_empty;
  wire _myaxi_write_req_fifo_almost_empty;

  _myaxi_write_req_fifo
  inst__myaxi_write_req_fifo
  (
    .CLK(CLK),
    .RST(RST),
    ._myaxi_write_req_fifo_enq(_myaxi_write_req_fifo_enq),
    ._myaxi_write_req_fifo_wdata(_myaxi_write_req_fifo_wdata),
    ._myaxi_write_req_fifo_full(_myaxi_write_req_fifo_full),
    ._myaxi_write_req_fifo_almost_full(_myaxi_write_req_fifo_almost_full),
    ._myaxi_write_req_fifo_deq(_myaxi_write_req_fifo_deq),
    ._myaxi_write_req_fifo_rdata(_myaxi_write_req_fifo_rdata),
    ._myaxi_write_req_fifo_empty(_myaxi_write_req_fifo_empty),
    ._myaxi_write_req_fifo_almost_empty(_myaxi_write_req_fifo_almost_empty)
  );

  reg [4-1:0] count__myaxi_write_req_fifo;
  wire [8-1:0] _myaxi_write_op_sel_fifo;
  wire [32-1:0] _myaxi_write_local_addr_fifo;
  wire [32-1:0] _myaxi_write_local_stride_fifo;
  wire [33-1:0] _myaxi_write_size_fifo;
  wire [32-1:0] _myaxi_write_local_blocksize_fifo;
  wire [8-1:0] unpack_write_req_op_sel_6;
  wire [32-1:0] unpack_write_req_local_addr_7;
  wire [32-1:0] unpack_write_req_local_stride_8;
  wire [33-1:0] unpack_write_req_size_9;
  wire [32-1:0] unpack_write_req_local_blocksize_10;
  assign unpack_write_req_op_sel_6 = _myaxi_write_req_fifo_rdata[136:129];
  assign unpack_write_req_local_addr_7 = _myaxi_write_req_fifo_rdata[128:97];
  assign unpack_write_req_local_stride_8 = _myaxi_write_req_fifo_rdata[96:65];
  assign unpack_write_req_size_9 = _myaxi_write_req_fifo_rdata[64:32];
  assign unpack_write_req_local_blocksize_10 = _myaxi_write_req_fifo_rdata[31:0];
  assign _myaxi_write_op_sel_fifo = unpack_write_req_op_sel_6;
  assign _myaxi_write_local_addr_fifo = unpack_write_req_local_addr_7;
  assign _myaxi_write_local_stride_fifo = unpack_write_req_local_stride_8;
  assign _myaxi_write_size_fifo = unpack_write_req_size_9;
  assign _myaxi_write_local_blocksize_fifo = unpack_write_req_local_blocksize_10;
  reg [8-1:0] _myaxi_write_op_sel_buf;
  reg [32-1:0] _myaxi_write_local_addr_buf;
  reg [32-1:0] _myaxi_write_local_stride_buf;
  reg [33-1:0] _myaxi_write_size_buf;
  reg [32-1:0] _myaxi_write_local_blocksize_buf;
  reg _myaxi_write_req_idle;
  reg _myaxi_write_data_idle;
  wire _myaxi_write_idle;
  assign _myaxi_write_idle = !_myaxi_write_start && _myaxi_write_req_idle && _myaxi_write_req_fifo_empty && _myaxi_write_data_idle;
  wire [20-1:0] ram_a_0_0_addr;
  wire [32-1:0] ram_a_0_0_rdata;
  wire [32-1:0] ram_a_0_0_wdata;
  wire ram_a_0_0_wenable;
  wire ram_a_0_0_enable;

  ram_a_0
  inst_ram_a_0
  (
    .CLK(CLK),
    .ram_a_0_0_addr(ram_a_0_0_addr),
    .ram_a_0_0_rdata(ram_a_0_0_rdata),
    .ram_a_0_0_wdata(ram_a_0_0_wdata),
    .ram_a_0_0_wenable(ram_a_0_0_wenable),
    .ram_a_0_0_enable(ram_a_0_0_enable)
  );

  wire [20-1:0] ram_a_1_0_addr;
  wire [32-1:0] ram_a_1_0_rdata;
  wire [32-1:0] ram_a_1_0_wdata;
  wire ram_a_1_0_wenable;
  wire ram_a_1_0_enable;

  ram_a_1
  inst_ram_a_1
  (
    .CLK(CLK),
    .ram_a_1_0_addr(ram_a_1_0_addr),
    .ram_a_1_0_rdata(ram_a_1_0_rdata),
    .ram_a_1_0_wdata(ram_a_1_0_wdata),
    .ram_a_1_0_wenable(ram_a_1_0_wenable),
    .ram_a_1_0_enable(ram_a_1_0_enable)
  );

  wire [20-1:0] ram_a_2_0_addr;
  wire [32-1:0] ram_a_2_0_rdata;
  wire [32-1:0] ram_a_2_0_wdata;
  wire ram_a_2_0_wenable;
  wire ram_a_2_0_enable;

  ram_a_2
  inst_ram_a_2
  (
    .CLK(CLK),
    .ram_a_2_0_addr(ram_a_2_0_addr),
    .ram_a_2_0_rdata(ram_a_2_0_rdata),
    .ram_a_2_0_wdata(ram_a_2_0_wdata),
    .ram_a_2_0_wenable(ram_a_2_0_wenable),
    .ram_a_2_0_enable(ram_a_2_0_enable)
  );

  wire [20-1:0] ram_a_3_0_addr;
  wire [32-1:0] ram_a_3_0_rdata;
  wire [32-1:0] ram_a_3_0_wdata;
  wire ram_a_3_0_wenable;
  wire ram_a_3_0_enable;

  ram_a_3
  inst_ram_a_3
  (
    .CLK(CLK),
    .ram_a_3_0_addr(ram_a_3_0_addr),
    .ram_a_3_0_rdata(ram_a_3_0_rdata),
    .ram_a_3_0_wdata(ram_a_3_0_wdata),
    .ram_a_3_0_wenable(ram_a_3_0_wenable),
    .ram_a_3_0_enable(ram_a_3_0_enable)
  );

  wire [20-1:0] ram_a_4_0_addr;
  wire [32-1:0] ram_a_4_0_rdata;
  wire [32-1:0] ram_a_4_0_wdata;
  wire ram_a_4_0_wenable;
  wire ram_a_4_0_enable;

  ram_a_4
  inst_ram_a_4
  (
    .CLK(CLK),
    .ram_a_4_0_addr(ram_a_4_0_addr),
    .ram_a_4_0_rdata(ram_a_4_0_rdata),
    .ram_a_4_0_wdata(ram_a_4_0_wdata),
    .ram_a_4_0_wenable(ram_a_4_0_wenable),
    .ram_a_4_0_enable(ram_a_4_0_enable)
  );

  wire [20-1:0] ram_a_5_0_addr;
  wire [32-1:0] ram_a_5_0_rdata;
  wire [32-1:0] ram_a_5_0_wdata;
  wire ram_a_5_0_wenable;
  wire ram_a_5_0_enable;

  ram_a_5
  inst_ram_a_5
  (
    .CLK(CLK),
    .ram_a_5_0_addr(ram_a_5_0_addr),
    .ram_a_5_0_rdata(ram_a_5_0_rdata),
    .ram_a_5_0_wdata(ram_a_5_0_wdata),
    .ram_a_5_0_wenable(ram_a_5_0_wenable),
    .ram_a_5_0_enable(ram_a_5_0_enable)
  );

  wire [20-1:0] ram_a_6_0_addr;
  wire [32-1:0] ram_a_6_0_rdata;
  wire [32-1:0] ram_a_6_0_wdata;
  wire ram_a_6_0_wenable;
  wire ram_a_6_0_enable;

  ram_a_6
  inst_ram_a_6
  (
    .CLK(CLK),
    .ram_a_6_0_addr(ram_a_6_0_addr),
    .ram_a_6_0_rdata(ram_a_6_0_rdata),
    .ram_a_6_0_wdata(ram_a_6_0_wdata),
    .ram_a_6_0_wenable(ram_a_6_0_wenable),
    .ram_a_6_0_enable(ram_a_6_0_enable)
  );

  wire [20-1:0] ram_a_7_0_addr;
  wire [32-1:0] ram_a_7_0_rdata;
  wire [32-1:0] ram_a_7_0_wdata;
  wire ram_a_7_0_wenable;
  wire ram_a_7_0_enable;

  ram_a_7
  inst_ram_a_7
  (
    .CLK(CLK),
    .ram_a_7_0_addr(ram_a_7_0_addr),
    .ram_a_7_0_rdata(ram_a_7_0_rdata),
    .ram_a_7_0_wdata(ram_a_7_0_wdata),
    .ram_a_7_0_wenable(ram_a_7_0_wenable),
    .ram_a_7_0_enable(ram_a_7_0_enable)
  );

  wire [20-1:0] ram_a_8_0_addr;
  wire [32-1:0] ram_a_8_0_rdata;
  wire [32-1:0] ram_a_8_0_wdata;
  wire ram_a_8_0_wenable;
  wire ram_a_8_0_enable;

  ram_a_8
  inst_ram_a_8
  (
    .CLK(CLK),
    .ram_a_8_0_addr(ram_a_8_0_addr),
    .ram_a_8_0_rdata(ram_a_8_0_rdata),
    .ram_a_8_0_wdata(ram_a_8_0_wdata),
    .ram_a_8_0_wenable(ram_a_8_0_wenable),
    .ram_a_8_0_enable(ram_a_8_0_enable)
  );

  wire [20-1:0] ram_a_9_0_addr;
  wire [32-1:0] ram_a_9_0_rdata;
  wire [32-1:0] ram_a_9_0_wdata;
  wire ram_a_9_0_wenable;
  wire ram_a_9_0_enable;

  ram_a_9
  inst_ram_a_9
  (
    .CLK(CLK),
    .ram_a_9_0_addr(ram_a_9_0_addr),
    .ram_a_9_0_rdata(ram_a_9_0_rdata),
    .ram_a_9_0_wdata(ram_a_9_0_wdata),
    .ram_a_9_0_wenable(ram_a_9_0_wenable),
    .ram_a_9_0_enable(ram_a_9_0_enable)
  );

  wire [20-1:0] ram_a_10_0_addr;
  wire [32-1:0] ram_a_10_0_rdata;
  wire [32-1:0] ram_a_10_0_wdata;
  wire ram_a_10_0_wenable;
  wire ram_a_10_0_enable;

  ram_a_10
  inst_ram_a_10
  (
    .CLK(CLK),
    .ram_a_10_0_addr(ram_a_10_0_addr),
    .ram_a_10_0_rdata(ram_a_10_0_rdata),
    .ram_a_10_0_wdata(ram_a_10_0_wdata),
    .ram_a_10_0_wenable(ram_a_10_0_wenable),
    .ram_a_10_0_enable(ram_a_10_0_enable)
  );

  wire [20-1:0] ram_a_11_0_addr;
  wire [32-1:0] ram_a_11_0_rdata;
  wire [32-1:0] ram_a_11_0_wdata;
  wire ram_a_11_0_wenable;
  wire ram_a_11_0_enable;

  ram_a_11
  inst_ram_a_11
  (
    .CLK(CLK),
    .ram_a_11_0_addr(ram_a_11_0_addr),
    .ram_a_11_0_rdata(ram_a_11_0_rdata),
    .ram_a_11_0_wdata(ram_a_11_0_wdata),
    .ram_a_11_0_wenable(ram_a_11_0_wenable),
    .ram_a_11_0_enable(ram_a_11_0_enable)
  );

  wire [20-1:0] ram_a_12_0_addr;
  wire [32-1:0] ram_a_12_0_rdata;
  wire [32-1:0] ram_a_12_0_wdata;
  wire ram_a_12_0_wenable;
  wire ram_a_12_0_enable;

  ram_a_12
  inst_ram_a_12
  (
    .CLK(CLK),
    .ram_a_12_0_addr(ram_a_12_0_addr),
    .ram_a_12_0_rdata(ram_a_12_0_rdata),
    .ram_a_12_0_wdata(ram_a_12_0_wdata),
    .ram_a_12_0_wenable(ram_a_12_0_wenable),
    .ram_a_12_0_enable(ram_a_12_0_enable)
  );

  wire [20-1:0] ram_a_13_0_addr;
  wire [32-1:0] ram_a_13_0_rdata;
  wire [32-1:0] ram_a_13_0_wdata;
  wire ram_a_13_0_wenable;
  wire ram_a_13_0_enable;

  ram_a_13
  inst_ram_a_13
  (
    .CLK(CLK),
    .ram_a_13_0_addr(ram_a_13_0_addr),
    .ram_a_13_0_rdata(ram_a_13_0_rdata),
    .ram_a_13_0_wdata(ram_a_13_0_wdata),
    .ram_a_13_0_wenable(ram_a_13_0_wenable),
    .ram_a_13_0_enable(ram_a_13_0_enable)
  );

  wire [20-1:0] ram_a_14_0_addr;
  wire [32-1:0] ram_a_14_0_rdata;
  wire [32-1:0] ram_a_14_0_wdata;
  wire ram_a_14_0_wenable;
  wire ram_a_14_0_enable;

  ram_a_14
  inst_ram_a_14
  (
    .CLK(CLK),
    .ram_a_14_0_addr(ram_a_14_0_addr),
    .ram_a_14_0_rdata(ram_a_14_0_rdata),
    .ram_a_14_0_wdata(ram_a_14_0_wdata),
    .ram_a_14_0_wenable(ram_a_14_0_wenable),
    .ram_a_14_0_enable(ram_a_14_0_enable)
  );

  wire [20-1:0] ram_a_15_0_addr;
  wire [32-1:0] ram_a_15_0_rdata;
  wire [32-1:0] ram_a_15_0_wdata;
  wire ram_a_15_0_wenable;
  wire ram_a_15_0_enable;

  ram_a_15
  inst_ram_a_15
  (
    .CLK(CLK),
    .ram_a_15_0_addr(ram_a_15_0_addr),
    .ram_a_15_0_rdata(ram_a_15_0_rdata),
    .ram_a_15_0_wdata(ram_a_15_0_wdata),
    .ram_a_15_0_wenable(ram_a_15_0_wenable),
    .ram_a_15_0_enable(ram_a_15_0_enable)
  );

  wire [20-1:0] ram_a_16_0_addr;
  wire [32-1:0] ram_a_16_0_rdata;
  wire [32-1:0] ram_a_16_0_wdata;
  wire ram_a_16_0_wenable;
  wire ram_a_16_0_enable;

  ram_a_16
  inst_ram_a_16
  (
    .CLK(CLK),
    .ram_a_16_0_addr(ram_a_16_0_addr),
    .ram_a_16_0_rdata(ram_a_16_0_rdata),
    .ram_a_16_0_wdata(ram_a_16_0_wdata),
    .ram_a_16_0_wenable(ram_a_16_0_wenable),
    .ram_a_16_0_enable(ram_a_16_0_enable)
  );

  wire [20-1:0] ram_a_17_0_addr;
  wire [32-1:0] ram_a_17_0_rdata;
  wire [32-1:0] ram_a_17_0_wdata;
  wire ram_a_17_0_wenable;
  wire ram_a_17_0_enable;

  ram_a_17
  inst_ram_a_17
  (
    .CLK(CLK),
    .ram_a_17_0_addr(ram_a_17_0_addr),
    .ram_a_17_0_rdata(ram_a_17_0_rdata),
    .ram_a_17_0_wdata(ram_a_17_0_wdata),
    .ram_a_17_0_wenable(ram_a_17_0_wenable),
    .ram_a_17_0_enable(ram_a_17_0_enable)
  );

  wire [20-1:0] ram_a_18_0_addr;
  wire [32-1:0] ram_a_18_0_rdata;
  wire [32-1:0] ram_a_18_0_wdata;
  wire ram_a_18_0_wenable;
  wire ram_a_18_0_enable;

  ram_a_18
  inst_ram_a_18
  (
    .CLK(CLK),
    .ram_a_18_0_addr(ram_a_18_0_addr),
    .ram_a_18_0_rdata(ram_a_18_0_rdata),
    .ram_a_18_0_wdata(ram_a_18_0_wdata),
    .ram_a_18_0_wenable(ram_a_18_0_wenable),
    .ram_a_18_0_enable(ram_a_18_0_enable)
  );

  wire [20-1:0] ram_a_19_0_addr;
  wire [32-1:0] ram_a_19_0_rdata;
  wire [32-1:0] ram_a_19_0_wdata;
  wire ram_a_19_0_wenable;
  wire ram_a_19_0_enable;

  ram_a_19
  inst_ram_a_19
  (
    .CLK(CLK),
    .ram_a_19_0_addr(ram_a_19_0_addr),
    .ram_a_19_0_rdata(ram_a_19_0_rdata),
    .ram_a_19_0_wdata(ram_a_19_0_wdata),
    .ram_a_19_0_wenable(ram_a_19_0_wenable),
    .ram_a_19_0_enable(ram_a_19_0_enable)
  );

  wire [20-1:0] ram_a_20_0_addr;
  wire [32-1:0] ram_a_20_0_rdata;
  wire [32-1:0] ram_a_20_0_wdata;
  wire ram_a_20_0_wenable;
  wire ram_a_20_0_enable;

  ram_a_20
  inst_ram_a_20
  (
    .CLK(CLK),
    .ram_a_20_0_addr(ram_a_20_0_addr),
    .ram_a_20_0_rdata(ram_a_20_0_rdata),
    .ram_a_20_0_wdata(ram_a_20_0_wdata),
    .ram_a_20_0_wenable(ram_a_20_0_wenable),
    .ram_a_20_0_enable(ram_a_20_0_enable)
  );

  wire [20-1:0] ram_a_21_0_addr;
  wire [32-1:0] ram_a_21_0_rdata;
  wire [32-1:0] ram_a_21_0_wdata;
  wire ram_a_21_0_wenable;
  wire ram_a_21_0_enable;

  ram_a_21
  inst_ram_a_21
  (
    .CLK(CLK),
    .ram_a_21_0_addr(ram_a_21_0_addr),
    .ram_a_21_0_rdata(ram_a_21_0_rdata),
    .ram_a_21_0_wdata(ram_a_21_0_wdata),
    .ram_a_21_0_wenable(ram_a_21_0_wenable),
    .ram_a_21_0_enable(ram_a_21_0_enable)
  );

  wire [20-1:0] ram_a_22_0_addr;
  wire [32-1:0] ram_a_22_0_rdata;
  wire [32-1:0] ram_a_22_0_wdata;
  wire ram_a_22_0_wenable;
  wire ram_a_22_0_enable;

  ram_a_22
  inst_ram_a_22
  (
    .CLK(CLK),
    .ram_a_22_0_addr(ram_a_22_0_addr),
    .ram_a_22_0_rdata(ram_a_22_0_rdata),
    .ram_a_22_0_wdata(ram_a_22_0_wdata),
    .ram_a_22_0_wenable(ram_a_22_0_wenable),
    .ram_a_22_0_enable(ram_a_22_0_enable)
  );

  wire [20-1:0] ram_a_23_0_addr;
  wire [32-1:0] ram_a_23_0_rdata;
  wire [32-1:0] ram_a_23_0_wdata;
  wire ram_a_23_0_wenable;
  wire ram_a_23_0_enable;

  ram_a_23
  inst_ram_a_23
  (
    .CLK(CLK),
    .ram_a_23_0_addr(ram_a_23_0_addr),
    .ram_a_23_0_rdata(ram_a_23_0_rdata),
    .ram_a_23_0_wdata(ram_a_23_0_wdata),
    .ram_a_23_0_wenable(ram_a_23_0_wenable),
    .ram_a_23_0_enable(ram_a_23_0_enable)
  );

  wire [20-1:0] ram_a_24_0_addr;
  wire [32-1:0] ram_a_24_0_rdata;
  wire [32-1:0] ram_a_24_0_wdata;
  wire ram_a_24_0_wenable;
  wire ram_a_24_0_enable;

  ram_a_24
  inst_ram_a_24
  (
    .CLK(CLK),
    .ram_a_24_0_addr(ram_a_24_0_addr),
    .ram_a_24_0_rdata(ram_a_24_0_rdata),
    .ram_a_24_0_wdata(ram_a_24_0_wdata),
    .ram_a_24_0_wenable(ram_a_24_0_wenable),
    .ram_a_24_0_enable(ram_a_24_0_enable)
  );

  wire [20-1:0] ram_a_25_0_addr;
  wire [32-1:0] ram_a_25_0_rdata;
  wire [32-1:0] ram_a_25_0_wdata;
  wire ram_a_25_0_wenable;
  wire ram_a_25_0_enable;

  ram_a_25
  inst_ram_a_25
  (
    .CLK(CLK),
    .ram_a_25_0_addr(ram_a_25_0_addr),
    .ram_a_25_0_rdata(ram_a_25_0_rdata),
    .ram_a_25_0_wdata(ram_a_25_0_wdata),
    .ram_a_25_0_wenable(ram_a_25_0_wenable),
    .ram_a_25_0_enable(ram_a_25_0_enable)
  );

  wire [20-1:0] ram_a_26_0_addr;
  wire [32-1:0] ram_a_26_0_rdata;
  wire [32-1:0] ram_a_26_0_wdata;
  wire ram_a_26_0_wenable;
  wire ram_a_26_0_enable;

  ram_a_26
  inst_ram_a_26
  (
    .CLK(CLK),
    .ram_a_26_0_addr(ram_a_26_0_addr),
    .ram_a_26_0_rdata(ram_a_26_0_rdata),
    .ram_a_26_0_wdata(ram_a_26_0_wdata),
    .ram_a_26_0_wenable(ram_a_26_0_wenable),
    .ram_a_26_0_enable(ram_a_26_0_enable)
  );

  wire [20-1:0] ram_a_27_0_addr;
  wire [32-1:0] ram_a_27_0_rdata;
  wire [32-1:0] ram_a_27_0_wdata;
  wire ram_a_27_0_wenable;
  wire ram_a_27_0_enable;

  ram_a_27
  inst_ram_a_27
  (
    .CLK(CLK),
    .ram_a_27_0_addr(ram_a_27_0_addr),
    .ram_a_27_0_rdata(ram_a_27_0_rdata),
    .ram_a_27_0_wdata(ram_a_27_0_wdata),
    .ram_a_27_0_wenable(ram_a_27_0_wenable),
    .ram_a_27_0_enable(ram_a_27_0_enable)
  );

  wire [20-1:0] ram_a_28_0_addr;
  wire [32-1:0] ram_a_28_0_rdata;
  wire [32-1:0] ram_a_28_0_wdata;
  wire ram_a_28_0_wenable;
  wire ram_a_28_0_enable;

  ram_a_28
  inst_ram_a_28
  (
    .CLK(CLK),
    .ram_a_28_0_addr(ram_a_28_0_addr),
    .ram_a_28_0_rdata(ram_a_28_0_rdata),
    .ram_a_28_0_wdata(ram_a_28_0_wdata),
    .ram_a_28_0_wenable(ram_a_28_0_wenable),
    .ram_a_28_0_enable(ram_a_28_0_enable)
  );

  wire [20-1:0] ram_a_29_0_addr;
  wire [32-1:0] ram_a_29_0_rdata;
  wire [32-1:0] ram_a_29_0_wdata;
  wire ram_a_29_0_wenable;
  wire ram_a_29_0_enable;

  ram_a_29
  inst_ram_a_29
  (
    .CLK(CLK),
    .ram_a_29_0_addr(ram_a_29_0_addr),
    .ram_a_29_0_rdata(ram_a_29_0_rdata),
    .ram_a_29_0_wdata(ram_a_29_0_wdata),
    .ram_a_29_0_wenable(ram_a_29_0_wenable),
    .ram_a_29_0_enable(ram_a_29_0_enable)
  );

  wire [20-1:0] ram_a_30_0_addr;
  wire [32-1:0] ram_a_30_0_rdata;
  wire [32-1:0] ram_a_30_0_wdata;
  wire ram_a_30_0_wenable;
  wire ram_a_30_0_enable;

  ram_a_30
  inst_ram_a_30
  (
    .CLK(CLK),
    .ram_a_30_0_addr(ram_a_30_0_addr),
    .ram_a_30_0_rdata(ram_a_30_0_rdata),
    .ram_a_30_0_wdata(ram_a_30_0_wdata),
    .ram_a_30_0_wenable(ram_a_30_0_wenable),
    .ram_a_30_0_enable(ram_a_30_0_enable)
  );

  wire [20-1:0] ram_a_31_0_addr;
  wire [32-1:0] ram_a_31_0_rdata;
  wire [32-1:0] ram_a_31_0_wdata;
  wire ram_a_31_0_wenable;
  wire ram_a_31_0_enable;

  ram_a_31
  inst_ram_a_31
  (
    .CLK(CLK),
    .ram_a_31_0_addr(ram_a_31_0_addr),
    .ram_a_31_0_rdata(ram_a_31_0_rdata),
    .ram_a_31_0_wdata(ram_a_31_0_wdata),
    .ram_a_31_0_wenable(ram_a_31_0_wenable),
    .ram_a_31_0_enable(ram_a_31_0_enable)
  );

  wire [20-1:0] ram_b_0_0_addr;
  wire [32-1:0] ram_b_0_0_rdata;
  wire [32-1:0] ram_b_0_0_wdata;
  wire ram_b_0_0_wenable;
  wire ram_b_0_0_enable;

  ram_b_0
  inst_ram_b_0
  (
    .CLK(CLK),
    .ram_b_0_0_addr(ram_b_0_0_addr),
    .ram_b_0_0_rdata(ram_b_0_0_rdata),
    .ram_b_0_0_wdata(ram_b_0_0_wdata),
    .ram_b_0_0_wenable(ram_b_0_0_wenable),
    .ram_b_0_0_enable(ram_b_0_0_enable)
  );

  wire [20-1:0] ram_b_1_0_addr;
  wire [32-1:0] ram_b_1_0_rdata;
  wire [32-1:0] ram_b_1_0_wdata;
  wire ram_b_1_0_wenable;
  wire ram_b_1_0_enable;

  ram_b_1
  inst_ram_b_1
  (
    .CLK(CLK),
    .ram_b_1_0_addr(ram_b_1_0_addr),
    .ram_b_1_0_rdata(ram_b_1_0_rdata),
    .ram_b_1_0_wdata(ram_b_1_0_wdata),
    .ram_b_1_0_wenable(ram_b_1_0_wenable),
    .ram_b_1_0_enable(ram_b_1_0_enable)
  );

  wire [20-1:0] ram_b_2_0_addr;
  wire [32-1:0] ram_b_2_0_rdata;
  wire [32-1:0] ram_b_2_0_wdata;
  wire ram_b_2_0_wenable;
  wire ram_b_2_0_enable;

  ram_b_2
  inst_ram_b_2
  (
    .CLK(CLK),
    .ram_b_2_0_addr(ram_b_2_0_addr),
    .ram_b_2_0_rdata(ram_b_2_0_rdata),
    .ram_b_2_0_wdata(ram_b_2_0_wdata),
    .ram_b_2_0_wenable(ram_b_2_0_wenable),
    .ram_b_2_0_enable(ram_b_2_0_enable)
  );

  wire [20-1:0] ram_b_3_0_addr;
  wire [32-1:0] ram_b_3_0_rdata;
  wire [32-1:0] ram_b_3_0_wdata;
  wire ram_b_3_0_wenable;
  wire ram_b_3_0_enable;

  ram_b_3
  inst_ram_b_3
  (
    .CLK(CLK),
    .ram_b_3_0_addr(ram_b_3_0_addr),
    .ram_b_3_0_rdata(ram_b_3_0_rdata),
    .ram_b_3_0_wdata(ram_b_3_0_wdata),
    .ram_b_3_0_wenable(ram_b_3_0_wenable),
    .ram_b_3_0_enable(ram_b_3_0_enable)
  );

  wire [20-1:0] ram_b_4_0_addr;
  wire [32-1:0] ram_b_4_0_rdata;
  wire [32-1:0] ram_b_4_0_wdata;
  wire ram_b_4_0_wenable;
  wire ram_b_4_0_enable;

  ram_b_4
  inst_ram_b_4
  (
    .CLK(CLK),
    .ram_b_4_0_addr(ram_b_4_0_addr),
    .ram_b_4_0_rdata(ram_b_4_0_rdata),
    .ram_b_4_0_wdata(ram_b_4_0_wdata),
    .ram_b_4_0_wenable(ram_b_4_0_wenable),
    .ram_b_4_0_enable(ram_b_4_0_enable)
  );

  wire [20-1:0] ram_b_5_0_addr;
  wire [32-1:0] ram_b_5_0_rdata;
  wire [32-1:0] ram_b_5_0_wdata;
  wire ram_b_5_0_wenable;
  wire ram_b_5_0_enable;

  ram_b_5
  inst_ram_b_5
  (
    .CLK(CLK),
    .ram_b_5_0_addr(ram_b_5_0_addr),
    .ram_b_5_0_rdata(ram_b_5_0_rdata),
    .ram_b_5_0_wdata(ram_b_5_0_wdata),
    .ram_b_5_0_wenable(ram_b_5_0_wenable),
    .ram_b_5_0_enable(ram_b_5_0_enable)
  );

  wire [20-1:0] ram_b_6_0_addr;
  wire [32-1:0] ram_b_6_0_rdata;
  wire [32-1:0] ram_b_6_0_wdata;
  wire ram_b_6_0_wenable;
  wire ram_b_6_0_enable;

  ram_b_6
  inst_ram_b_6
  (
    .CLK(CLK),
    .ram_b_6_0_addr(ram_b_6_0_addr),
    .ram_b_6_0_rdata(ram_b_6_0_rdata),
    .ram_b_6_0_wdata(ram_b_6_0_wdata),
    .ram_b_6_0_wenable(ram_b_6_0_wenable),
    .ram_b_6_0_enable(ram_b_6_0_enable)
  );

  wire [20-1:0] ram_b_7_0_addr;
  wire [32-1:0] ram_b_7_0_rdata;
  wire [32-1:0] ram_b_7_0_wdata;
  wire ram_b_7_0_wenable;
  wire ram_b_7_0_enable;

  ram_b_7
  inst_ram_b_7
  (
    .CLK(CLK),
    .ram_b_7_0_addr(ram_b_7_0_addr),
    .ram_b_7_0_rdata(ram_b_7_0_rdata),
    .ram_b_7_0_wdata(ram_b_7_0_wdata),
    .ram_b_7_0_wenable(ram_b_7_0_wenable),
    .ram_b_7_0_enable(ram_b_7_0_enable)
  );

  wire [20-1:0] ram_b_8_0_addr;
  wire [32-1:0] ram_b_8_0_rdata;
  wire [32-1:0] ram_b_8_0_wdata;
  wire ram_b_8_0_wenable;
  wire ram_b_8_0_enable;

  ram_b_8
  inst_ram_b_8
  (
    .CLK(CLK),
    .ram_b_8_0_addr(ram_b_8_0_addr),
    .ram_b_8_0_rdata(ram_b_8_0_rdata),
    .ram_b_8_0_wdata(ram_b_8_0_wdata),
    .ram_b_8_0_wenable(ram_b_8_0_wenable),
    .ram_b_8_0_enable(ram_b_8_0_enable)
  );

  wire [20-1:0] ram_b_9_0_addr;
  wire [32-1:0] ram_b_9_0_rdata;
  wire [32-1:0] ram_b_9_0_wdata;
  wire ram_b_9_0_wenable;
  wire ram_b_9_0_enable;

  ram_b_9
  inst_ram_b_9
  (
    .CLK(CLK),
    .ram_b_9_0_addr(ram_b_9_0_addr),
    .ram_b_9_0_rdata(ram_b_9_0_rdata),
    .ram_b_9_0_wdata(ram_b_9_0_wdata),
    .ram_b_9_0_wenable(ram_b_9_0_wenable),
    .ram_b_9_0_enable(ram_b_9_0_enable)
  );

  wire [20-1:0] ram_b_10_0_addr;
  wire [32-1:0] ram_b_10_0_rdata;
  wire [32-1:0] ram_b_10_0_wdata;
  wire ram_b_10_0_wenable;
  wire ram_b_10_0_enable;

  ram_b_10
  inst_ram_b_10
  (
    .CLK(CLK),
    .ram_b_10_0_addr(ram_b_10_0_addr),
    .ram_b_10_0_rdata(ram_b_10_0_rdata),
    .ram_b_10_0_wdata(ram_b_10_0_wdata),
    .ram_b_10_0_wenable(ram_b_10_0_wenable),
    .ram_b_10_0_enable(ram_b_10_0_enable)
  );

  wire [20-1:0] ram_b_11_0_addr;
  wire [32-1:0] ram_b_11_0_rdata;
  wire [32-1:0] ram_b_11_0_wdata;
  wire ram_b_11_0_wenable;
  wire ram_b_11_0_enable;

  ram_b_11
  inst_ram_b_11
  (
    .CLK(CLK),
    .ram_b_11_0_addr(ram_b_11_0_addr),
    .ram_b_11_0_rdata(ram_b_11_0_rdata),
    .ram_b_11_0_wdata(ram_b_11_0_wdata),
    .ram_b_11_0_wenable(ram_b_11_0_wenable),
    .ram_b_11_0_enable(ram_b_11_0_enable)
  );

  wire [20-1:0] ram_b_12_0_addr;
  wire [32-1:0] ram_b_12_0_rdata;
  wire [32-1:0] ram_b_12_0_wdata;
  wire ram_b_12_0_wenable;
  wire ram_b_12_0_enable;

  ram_b_12
  inst_ram_b_12
  (
    .CLK(CLK),
    .ram_b_12_0_addr(ram_b_12_0_addr),
    .ram_b_12_0_rdata(ram_b_12_0_rdata),
    .ram_b_12_0_wdata(ram_b_12_0_wdata),
    .ram_b_12_0_wenable(ram_b_12_0_wenable),
    .ram_b_12_0_enable(ram_b_12_0_enable)
  );

  wire [20-1:0] ram_b_13_0_addr;
  wire [32-1:0] ram_b_13_0_rdata;
  wire [32-1:0] ram_b_13_0_wdata;
  wire ram_b_13_0_wenable;
  wire ram_b_13_0_enable;

  ram_b_13
  inst_ram_b_13
  (
    .CLK(CLK),
    .ram_b_13_0_addr(ram_b_13_0_addr),
    .ram_b_13_0_rdata(ram_b_13_0_rdata),
    .ram_b_13_0_wdata(ram_b_13_0_wdata),
    .ram_b_13_0_wenable(ram_b_13_0_wenable),
    .ram_b_13_0_enable(ram_b_13_0_enable)
  );

  wire [20-1:0] ram_b_14_0_addr;
  wire [32-1:0] ram_b_14_0_rdata;
  wire [32-1:0] ram_b_14_0_wdata;
  wire ram_b_14_0_wenable;
  wire ram_b_14_0_enable;

  ram_b_14
  inst_ram_b_14
  (
    .CLK(CLK),
    .ram_b_14_0_addr(ram_b_14_0_addr),
    .ram_b_14_0_rdata(ram_b_14_0_rdata),
    .ram_b_14_0_wdata(ram_b_14_0_wdata),
    .ram_b_14_0_wenable(ram_b_14_0_wenable),
    .ram_b_14_0_enable(ram_b_14_0_enable)
  );

  wire [20-1:0] ram_b_15_0_addr;
  wire [32-1:0] ram_b_15_0_rdata;
  wire [32-1:0] ram_b_15_0_wdata;
  wire ram_b_15_0_wenable;
  wire ram_b_15_0_enable;

  ram_b_15
  inst_ram_b_15
  (
    .CLK(CLK),
    .ram_b_15_0_addr(ram_b_15_0_addr),
    .ram_b_15_0_rdata(ram_b_15_0_rdata),
    .ram_b_15_0_wdata(ram_b_15_0_wdata),
    .ram_b_15_0_wenable(ram_b_15_0_wenable),
    .ram_b_15_0_enable(ram_b_15_0_enable)
  );

  wire [20-1:0] ram_b_16_0_addr;
  wire [32-1:0] ram_b_16_0_rdata;
  wire [32-1:0] ram_b_16_0_wdata;
  wire ram_b_16_0_wenable;
  wire ram_b_16_0_enable;

  ram_b_16
  inst_ram_b_16
  (
    .CLK(CLK),
    .ram_b_16_0_addr(ram_b_16_0_addr),
    .ram_b_16_0_rdata(ram_b_16_0_rdata),
    .ram_b_16_0_wdata(ram_b_16_0_wdata),
    .ram_b_16_0_wenable(ram_b_16_0_wenable),
    .ram_b_16_0_enable(ram_b_16_0_enable)
  );

  wire [20-1:0] ram_b_17_0_addr;
  wire [32-1:0] ram_b_17_0_rdata;
  wire [32-1:0] ram_b_17_0_wdata;
  wire ram_b_17_0_wenable;
  wire ram_b_17_0_enable;

  ram_b_17
  inst_ram_b_17
  (
    .CLK(CLK),
    .ram_b_17_0_addr(ram_b_17_0_addr),
    .ram_b_17_0_rdata(ram_b_17_0_rdata),
    .ram_b_17_0_wdata(ram_b_17_0_wdata),
    .ram_b_17_0_wenable(ram_b_17_0_wenable),
    .ram_b_17_0_enable(ram_b_17_0_enable)
  );

  wire [20-1:0] ram_b_18_0_addr;
  wire [32-1:0] ram_b_18_0_rdata;
  wire [32-1:0] ram_b_18_0_wdata;
  wire ram_b_18_0_wenable;
  wire ram_b_18_0_enable;

  ram_b_18
  inst_ram_b_18
  (
    .CLK(CLK),
    .ram_b_18_0_addr(ram_b_18_0_addr),
    .ram_b_18_0_rdata(ram_b_18_0_rdata),
    .ram_b_18_0_wdata(ram_b_18_0_wdata),
    .ram_b_18_0_wenable(ram_b_18_0_wenable),
    .ram_b_18_0_enable(ram_b_18_0_enable)
  );

  wire [20-1:0] ram_b_19_0_addr;
  wire [32-1:0] ram_b_19_0_rdata;
  wire [32-1:0] ram_b_19_0_wdata;
  wire ram_b_19_0_wenable;
  wire ram_b_19_0_enable;

  ram_b_19
  inst_ram_b_19
  (
    .CLK(CLK),
    .ram_b_19_0_addr(ram_b_19_0_addr),
    .ram_b_19_0_rdata(ram_b_19_0_rdata),
    .ram_b_19_0_wdata(ram_b_19_0_wdata),
    .ram_b_19_0_wenable(ram_b_19_0_wenable),
    .ram_b_19_0_enable(ram_b_19_0_enable)
  );

  wire [20-1:0] ram_b_20_0_addr;
  wire [32-1:0] ram_b_20_0_rdata;
  wire [32-1:0] ram_b_20_0_wdata;
  wire ram_b_20_0_wenable;
  wire ram_b_20_0_enable;

  ram_b_20
  inst_ram_b_20
  (
    .CLK(CLK),
    .ram_b_20_0_addr(ram_b_20_0_addr),
    .ram_b_20_0_rdata(ram_b_20_0_rdata),
    .ram_b_20_0_wdata(ram_b_20_0_wdata),
    .ram_b_20_0_wenable(ram_b_20_0_wenable),
    .ram_b_20_0_enable(ram_b_20_0_enable)
  );

  wire [20-1:0] ram_b_21_0_addr;
  wire [32-1:0] ram_b_21_0_rdata;
  wire [32-1:0] ram_b_21_0_wdata;
  wire ram_b_21_0_wenable;
  wire ram_b_21_0_enable;

  ram_b_21
  inst_ram_b_21
  (
    .CLK(CLK),
    .ram_b_21_0_addr(ram_b_21_0_addr),
    .ram_b_21_0_rdata(ram_b_21_0_rdata),
    .ram_b_21_0_wdata(ram_b_21_0_wdata),
    .ram_b_21_0_wenable(ram_b_21_0_wenable),
    .ram_b_21_0_enable(ram_b_21_0_enable)
  );

  wire [20-1:0] ram_b_22_0_addr;
  wire [32-1:0] ram_b_22_0_rdata;
  wire [32-1:0] ram_b_22_0_wdata;
  wire ram_b_22_0_wenable;
  wire ram_b_22_0_enable;

  ram_b_22
  inst_ram_b_22
  (
    .CLK(CLK),
    .ram_b_22_0_addr(ram_b_22_0_addr),
    .ram_b_22_0_rdata(ram_b_22_0_rdata),
    .ram_b_22_0_wdata(ram_b_22_0_wdata),
    .ram_b_22_0_wenable(ram_b_22_0_wenable),
    .ram_b_22_0_enable(ram_b_22_0_enable)
  );

  wire [20-1:0] ram_b_23_0_addr;
  wire [32-1:0] ram_b_23_0_rdata;
  wire [32-1:0] ram_b_23_0_wdata;
  wire ram_b_23_0_wenable;
  wire ram_b_23_0_enable;

  ram_b_23
  inst_ram_b_23
  (
    .CLK(CLK),
    .ram_b_23_0_addr(ram_b_23_0_addr),
    .ram_b_23_0_rdata(ram_b_23_0_rdata),
    .ram_b_23_0_wdata(ram_b_23_0_wdata),
    .ram_b_23_0_wenable(ram_b_23_0_wenable),
    .ram_b_23_0_enable(ram_b_23_0_enable)
  );

  wire [20-1:0] ram_b_24_0_addr;
  wire [32-1:0] ram_b_24_0_rdata;
  wire [32-1:0] ram_b_24_0_wdata;
  wire ram_b_24_0_wenable;
  wire ram_b_24_0_enable;

  ram_b_24
  inst_ram_b_24
  (
    .CLK(CLK),
    .ram_b_24_0_addr(ram_b_24_0_addr),
    .ram_b_24_0_rdata(ram_b_24_0_rdata),
    .ram_b_24_0_wdata(ram_b_24_0_wdata),
    .ram_b_24_0_wenable(ram_b_24_0_wenable),
    .ram_b_24_0_enable(ram_b_24_0_enable)
  );

  wire [20-1:0] ram_b_25_0_addr;
  wire [32-1:0] ram_b_25_0_rdata;
  wire [32-1:0] ram_b_25_0_wdata;
  wire ram_b_25_0_wenable;
  wire ram_b_25_0_enable;

  ram_b_25
  inst_ram_b_25
  (
    .CLK(CLK),
    .ram_b_25_0_addr(ram_b_25_0_addr),
    .ram_b_25_0_rdata(ram_b_25_0_rdata),
    .ram_b_25_0_wdata(ram_b_25_0_wdata),
    .ram_b_25_0_wenable(ram_b_25_0_wenable),
    .ram_b_25_0_enable(ram_b_25_0_enable)
  );

  wire [20-1:0] ram_b_26_0_addr;
  wire [32-1:0] ram_b_26_0_rdata;
  wire [32-1:0] ram_b_26_0_wdata;
  wire ram_b_26_0_wenable;
  wire ram_b_26_0_enable;

  ram_b_26
  inst_ram_b_26
  (
    .CLK(CLK),
    .ram_b_26_0_addr(ram_b_26_0_addr),
    .ram_b_26_0_rdata(ram_b_26_0_rdata),
    .ram_b_26_0_wdata(ram_b_26_0_wdata),
    .ram_b_26_0_wenable(ram_b_26_0_wenable),
    .ram_b_26_0_enable(ram_b_26_0_enable)
  );

  wire [20-1:0] ram_b_27_0_addr;
  wire [32-1:0] ram_b_27_0_rdata;
  wire [32-1:0] ram_b_27_0_wdata;
  wire ram_b_27_0_wenable;
  wire ram_b_27_0_enable;

  ram_b_27
  inst_ram_b_27
  (
    .CLK(CLK),
    .ram_b_27_0_addr(ram_b_27_0_addr),
    .ram_b_27_0_rdata(ram_b_27_0_rdata),
    .ram_b_27_0_wdata(ram_b_27_0_wdata),
    .ram_b_27_0_wenable(ram_b_27_0_wenable),
    .ram_b_27_0_enable(ram_b_27_0_enable)
  );

  wire [20-1:0] ram_b_28_0_addr;
  wire [32-1:0] ram_b_28_0_rdata;
  wire [32-1:0] ram_b_28_0_wdata;
  wire ram_b_28_0_wenable;
  wire ram_b_28_0_enable;

  ram_b_28
  inst_ram_b_28
  (
    .CLK(CLK),
    .ram_b_28_0_addr(ram_b_28_0_addr),
    .ram_b_28_0_rdata(ram_b_28_0_rdata),
    .ram_b_28_0_wdata(ram_b_28_0_wdata),
    .ram_b_28_0_wenable(ram_b_28_0_wenable),
    .ram_b_28_0_enable(ram_b_28_0_enable)
  );

  wire [20-1:0] ram_b_29_0_addr;
  wire [32-1:0] ram_b_29_0_rdata;
  wire [32-1:0] ram_b_29_0_wdata;
  wire ram_b_29_0_wenable;
  wire ram_b_29_0_enable;

  ram_b_29
  inst_ram_b_29
  (
    .CLK(CLK),
    .ram_b_29_0_addr(ram_b_29_0_addr),
    .ram_b_29_0_rdata(ram_b_29_0_rdata),
    .ram_b_29_0_wdata(ram_b_29_0_wdata),
    .ram_b_29_0_wenable(ram_b_29_0_wenable),
    .ram_b_29_0_enable(ram_b_29_0_enable)
  );

  wire [20-1:0] ram_b_30_0_addr;
  wire [32-1:0] ram_b_30_0_rdata;
  wire [32-1:0] ram_b_30_0_wdata;
  wire ram_b_30_0_wenable;
  wire ram_b_30_0_enable;

  ram_b_30
  inst_ram_b_30
  (
    .CLK(CLK),
    .ram_b_30_0_addr(ram_b_30_0_addr),
    .ram_b_30_0_rdata(ram_b_30_0_rdata),
    .ram_b_30_0_wdata(ram_b_30_0_wdata),
    .ram_b_30_0_wenable(ram_b_30_0_wenable),
    .ram_b_30_0_enable(ram_b_30_0_enable)
  );

  wire [20-1:0] ram_b_31_0_addr;
  wire [32-1:0] ram_b_31_0_rdata;
  wire [32-1:0] ram_b_31_0_wdata;
  wire ram_b_31_0_wenable;
  wire ram_b_31_0_enable;

  ram_b_31
  inst_ram_b_31
  (
    .CLK(CLK),
    .ram_b_31_0_addr(ram_b_31_0_addr),
    .ram_b_31_0_rdata(ram_b_31_0_rdata),
    .ram_b_31_0_wdata(ram_b_31_0_wdata),
    .ram_b_31_0_wenable(ram_b_31_0_wenable),
    .ram_b_31_0_enable(ram_b_31_0_enable)
  );

  wire [20-1:0] ram_c_0_0_addr;
  wire [32-1:0] ram_c_0_0_rdata;
  wire [32-1:0] ram_c_0_0_wdata;
  wire ram_c_0_0_wenable;
  wire ram_c_0_0_enable;

  ram_c_0
  inst_ram_c_0
  (
    .CLK(CLK),
    .ram_c_0_0_addr(ram_c_0_0_addr),
    .ram_c_0_0_rdata(ram_c_0_0_rdata),
    .ram_c_0_0_wdata(ram_c_0_0_wdata),
    .ram_c_0_0_wenable(ram_c_0_0_wenable),
    .ram_c_0_0_enable(ram_c_0_0_enable)
  );

  wire [20-1:0] ram_c_1_0_addr;
  wire [32-1:0] ram_c_1_0_rdata;
  wire [32-1:0] ram_c_1_0_wdata;
  wire ram_c_1_0_wenable;
  wire ram_c_1_0_enable;

  ram_c_1
  inst_ram_c_1
  (
    .CLK(CLK),
    .ram_c_1_0_addr(ram_c_1_0_addr),
    .ram_c_1_0_rdata(ram_c_1_0_rdata),
    .ram_c_1_0_wdata(ram_c_1_0_wdata),
    .ram_c_1_0_wenable(ram_c_1_0_wenable),
    .ram_c_1_0_enable(ram_c_1_0_enable)
  );

  wire [20-1:0] ram_c_2_0_addr;
  wire [32-1:0] ram_c_2_0_rdata;
  wire [32-1:0] ram_c_2_0_wdata;
  wire ram_c_2_0_wenable;
  wire ram_c_2_0_enable;

  ram_c_2
  inst_ram_c_2
  (
    .CLK(CLK),
    .ram_c_2_0_addr(ram_c_2_0_addr),
    .ram_c_2_0_rdata(ram_c_2_0_rdata),
    .ram_c_2_0_wdata(ram_c_2_0_wdata),
    .ram_c_2_0_wenable(ram_c_2_0_wenable),
    .ram_c_2_0_enable(ram_c_2_0_enable)
  );

  wire [20-1:0] ram_c_3_0_addr;
  wire [32-1:0] ram_c_3_0_rdata;
  wire [32-1:0] ram_c_3_0_wdata;
  wire ram_c_3_0_wenable;
  wire ram_c_3_0_enable;

  ram_c_3
  inst_ram_c_3
  (
    .CLK(CLK),
    .ram_c_3_0_addr(ram_c_3_0_addr),
    .ram_c_3_0_rdata(ram_c_3_0_rdata),
    .ram_c_3_0_wdata(ram_c_3_0_wdata),
    .ram_c_3_0_wenable(ram_c_3_0_wenable),
    .ram_c_3_0_enable(ram_c_3_0_enable)
  );

  wire [20-1:0] ram_c_4_0_addr;
  wire [32-1:0] ram_c_4_0_rdata;
  wire [32-1:0] ram_c_4_0_wdata;
  wire ram_c_4_0_wenable;
  wire ram_c_4_0_enable;

  ram_c_4
  inst_ram_c_4
  (
    .CLK(CLK),
    .ram_c_4_0_addr(ram_c_4_0_addr),
    .ram_c_4_0_rdata(ram_c_4_0_rdata),
    .ram_c_4_0_wdata(ram_c_4_0_wdata),
    .ram_c_4_0_wenable(ram_c_4_0_wenable),
    .ram_c_4_0_enable(ram_c_4_0_enable)
  );

  wire [20-1:0] ram_c_5_0_addr;
  wire [32-1:0] ram_c_5_0_rdata;
  wire [32-1:0] ram_c_5_0_wdata;
  wire ram_c_5_0_wenable;
  wire ram_c_5_0_enable;

  ram_c_5
  inst_ram_c_5
  (
    .CLK(CLK),
    .ram_c_5_0_addr(ram_c_5_0_addr),
    .ram_c_5_0_rdata(ram_c_5_0_rdata),
    .ram_c_5_0_wdata(ram_c_5_0_wdata),
    .ram_c_5_0_wenable(ram_c_5_0_wenable),
    .ram_c_5_0_enable(ram_c_5_0_enable)
  );

  wire [20-1:0] ram_c_6_0_addr;
  wire [32-1:0] ram_c_6_0_rdata;
  wire [32-1:0] ram_c_6_0_wdata;
  wire ram_c_6_0_wenable;
  wire ram_c_6_0_enable;

  ram_c_6
  inst_ram_c_6
  (
    .CLK(CLK),
    .ram_c_6_0_addr(ram_c_6_0_addr),
    .ram_c_6_0_rdata(ram_c_6_0_rdata),
    .ram_c_6_0_wdata(ram_c_6_0_wdata),
    .ram_c_6_0_wenable(ram_c_6_0_wenable),
    .ram_c_6_0_enable(ram_c_6_0_enable)
  );

  wire [20-1:0] ram_c_7_0_addr;
  wire [32-1:0] ram_c_7_0_rdata;
  wire [32-1:0] ram_c_7_0_wdata;
  wire ram_c_7_0_wenable;
  wire ram_c_7_0_enable;

  ram_c_7
  inst_ram_c_7
  (
    .CLK(CLK),
    .ram_c_7_0_addr(ram_c_7_0_addr),
    .ram_c_7_0_rdata(ram_c_7_0_rdata),
    .ram_c_7_0_wdata(ram_c_7_0_wdata),
    .ram_c_7_0_wenable(ram_c_7_0_wenable),
    .ram_c_7_0_enable(ram_c_7_0_enable)
  );

  wire [20-1:0] ram_c_8_0_addr;
  wire [32-1:0] ram_c_8_0_rdata;
  wire [32-1:0] ram_c_8_0_wdata;
  wire ram_c_8_0_wenable;
  wire ram_c_8_0_enable;

  ram_c_8
  inst_ram_c_8
  (
    .CLK(CLK),
    .ram_c_8_0_addr(ram_c_8_0_addr),
    .ram_c_8_0_rdata(ram_c_8_0_rdata),
    .ram_c_8_0_wdata(ram_c_8_0_wdata),
    .ram_c_8_0_wenable(ram_c_8_0_wenable),
    .ram_c_8_0_enable(ram_c_8_0_enable)
  );

  wire [20-1:0] ram_c_9_0_addr;
  wire [32-1:0] ram_c_9_0_rdata;
  wire [32-1:0] ram_c_9_0_wdata;
  wire ram_c_9_0_wenable;
  wire ram_c_9_0_enable;

  ram_c_9
  inst_ram_c_9
  (
    .CLK(CLK),
    .ram_c_9_0_addr(ram_c_9_0_addr),
    .ram_c_9_0_rdata(ram_c_9_0_rdata),
    .ram_c_9_0_wdata(ram_c_9_0_wdata),
    .ram_c_9_0_wenable(ram_c_9_0_wenable),
    .ram_c_9_0_enable(ram_c_9_0_enable)
  );

  wire [20-1:0] ram_c_10_0_addr;
  wire [32-1:0] ram_c_10_0_rdata;
  wire [32-1:0] ram_c_10_0_wdata;
  wire ram_c_10_0_wenable;
  wire ram_c_10_0_enable;

  ram_c_10
  inst_ram_c_10
  (
    .CLK(CLK),
    .ram_c_10_0_addr(ram_c_10_0_addr),
    .ram_c_10_0_rdata(ram_c_10_0_rdata),
    .ram_c_10_0_wdata(ram_c_10_0_wdata),
    .ram_c_10_0_wenable(ram_c_10_0_wenable),
    .ram_c_10_0_enable(ram_c_10_0_enable)
  );

  wire [20-1:0] ram_c_11_0_addr;
  wire [32-1:0] ram_c_11_0_rdata;
  wire [32-1:0] ram_c_11_0_wdata;
  wire ram_c_11_0_wenable;
  wire ram_c_11_0_enable;

  ram_c_11
  inst_ram_c_11
  (
    .CLK(CLK),
    .ram_c_11_0_addr(ram_c_11_0_addr),
    .ram_c_11_0_rdata(ram_c_11_0_rdata),
    .ram_c_11_0_wdata(ram_c_11_0_wdata),
    .ram_c_11_0_wenable(ram_c_11_0_wenable),
    .ram_c_11_0_enable(ram_c_11_0_enable)
  );

  wire [20-1:0] ram_c_12_0_addr;
  wire [32-1:0] ram_c_12_0_rdata;
  wire [32-1:0] ram_c_12_0_wdata;
  wire ram_c_12_0_wenable;
  wire ram_c_12_0_enable;

  ram_c_12
  inst_ram_c_12
  (
    .CLK(CLK),
    .ram_c_12_0_addr(ram_c_12_0_addr),
    .ram_c_12_0_rdata(ram_c_12_0_rdata),
    .ram_c_12_0_wdata(ram_c_12_0_wdata),
    .ram_c_12_0_wenable(ram_c_12_0_wenable),
    .ram_c_12_0_enable(ram_c_12_0_enable)
  );

  wire [20-1:0] ram_c_13_0_addr;
  wire [32-1:0] ram_c_13_0_rdata;
  wire [32-1:0] ram_c_13_0_wdata;
  wire ram_c_13_0_wenable;
  wire ram_c_13_0_enable;

  ram_c_13
  inst_ram_c_13
  (
    .CLK(CLK),
    .ram_c_13_0_addr(ram_c_13_0_addr),
    .ram_c_13_0_rdata(ram_c_13_0_rdata),
    .ram_c_13_0_wdata(ram_c_13_0_wdata),
    .ram_c_13_0_wenable(ram_c_13_0_wenable),
    .ram_c_13_0_enable(ram_c_13_0_enable)
  );

  wire [20-1:0] ram_c_14_0_addr;
  wire [32-1:0] ram_c_14_0_rdata;
  wire [32-1:0] ram_c_14_0_wdata;
  wire ram_c_14_0_wenable;
  wire ram_c_14_0_enable;

  ram_c_14
  inst_ram_c_14
  (
    .CLK(CLK),
    .ram_c_14_0_addr(ram_c_14_0_addr),
    .ram_c_14_0_rdata(ram_c_14_0_rdata),
    .ram_c_14_0_wdata(ram_c_14_0_wdata),
    .ram_c_14_0_wenable(ram_c_14_0_wenable),
    .ram_c_14_0_enable(ram_c_14_0_enable)
  );

  wire [20-1:0] ram_c_15_0_addr;
  wire [32-1:0] ram_c_15_0_rdata;
  wire [32-1:0] ram_c_15_0_wdata;
  wire ram_c_15_0_wenable;
  wire ram_c_15_0_enable;

  ram_c_15
  inst_ram_c_15
  (
    .CLK(CLK),
    .ram_c_15_0_addr(ram_c_15_0_addr),
    .ram_c_15_0_rdata(ram_c_15_0_rdata),
    .ram_c_15_0_wdata(ram_c_15_0_wdata),
    .ram_c_15_0_wenable(ram_c_15_0_wenable),
    .ram_c_15_0_enable(ram_c_15_0_enable)
  );

  wire [20-1:0] ram_c_16_0_addr;
  wire [32-1:0] ram_c_16_0_rdata;
  wire [32-1:0] ram_c_16_0_wdata;
  wire ram_c_16_0_wenable;
  wire ram_c_16_0_enable;

  ram_c_16
  inst_ram_c_16
  (
    .CLK(CLK),
    .ram_c_16_0_addr(ram_c_16_0_addr),
    .ram_c_16_0_rdata(ram_c_16_0_rdata),
    .ram_c_16_0_wdata(ram_c_16_0_wdata),
    .ram_c_16_0_wenable(ram_c_16_0_wenable),
    .ram_c_16_0_enable(ram_c_16_0_enable)
  );

  wire [20-1:0] ram_c_17_0_addr;
  wire [32-1:0] ram_c_17_0_rdata;
  wire [32-1:0] ram_c_17_0_wdata;
  wire ram_c_17_0_wenable;
  wire ram_c_17_0_enable;

  ram_c_17
  inst_ram_c_17
  (
    .CLK(CLK),
    .ram_c_17_0_addr(ram_c_17_0_addr),
    .ram_c_17_0_rdata(ram_c_17_0_rdata),
    .ram_c_17_0_wdata(ram_c_17_0_wdata),
    .ram_c_17_0_wenable(ram_c_17_0_wenable),
    .ram_c_17_0_enable(ram_c_17_0_enable)
  );

  wire [20-1:0] ram_c_18_0_addr;
  wire [32-1:0] ram_c_18_0_rdata;
  wire [32-1:0] ram_c_18_0_wdata;
  wire ram_c_18_0_wenable;
  wire ram_c_18_0_enable;

  ram_c_18
  inst_ram_c_18
  (
    .CLK(CLK),
    .ram_c_18_0_addr(ram_c_18_0_addr),
    .ram_c_18_0_rdata(ram_c_18_0_rdata),
    .ram_c_18_0_wdata(ram_c_18_0_wdata),
    .ram_c_18_0_wenable(ram_c_18_0_wenable),
    .ram_c_18_0_enable(ram_c_18_0_enable)
  );

  wire [20-1:0] ram_c_19_0_addr;
  wire [32-1:0] ram_c_19_0_rdata;
  wire [32-1:0] ram_c_19_0_wdata;
  wire ram_c_19_0_wenable;
  wire ram_c_19_0_enable;

  ram_c_19
  inst_ram_c_19
  (
    .CLK(CLK),
    .ram_c_19_0_addr(ram_c_19_0_addr),
    .ram_c_19_0_rdata(ram_c_19_0_rdata),
    .ram_c_19_0_wdata(ram_c_19_0_wdata),
    .ram_c_19_0_wenable(ram_c_19_0_wenable),
    .ram_c_19_0_enable(ram_c_19_0_enable)
  );

  wire [20-1:0] ram_c_20_0_addr;
  wire [32-1:0] ram_c_20_0_rdata;
  wire [32-1:0] ram_c_20_0_wdata;
  wire ram_c_20_0_wenable;
  wire ram_c_20_0_enable;

  ram_c_20
  inst_ram_c_20
  (
    .CLK(CLK),
    .ram_c_20_0_addr(ram_c_20_0_addr),
    .ram_c_20_0_rdata(ram_c_20_0_rdata),
    .ram_c_20_0_wdata(ram_c_20_0_wdata),
    .ram_c_20_0_wenable(ram_c_20_0_wenable),
    .ram_c_20_0_enable(ram_c_20_0_enable)
  );

  wire [20-1:0] ram_c_21_0_addr;
  wire [32-1:0] ram_c_21_0_rdata;
  wire [32-1:0] ram_c_21_0_wdata;
  wire ram_c_21_0_wenable;
  wire ram_c_21_0_enable;

  ram_c_21
  inst_ram_c_21
  (
    .CLK(CLK),
    .ram_c_21_0_addr(ram_c_21_0_addr),
    .ram_c_21_0_rdata(ram_c_21_0_rdata),
    .ram_c_21_0_wdata(ram_c_21_0_wdata),
    .ram_c_21_0_wenable(ram_c_21_0_wenable),
    .ram_c_21_0_enable(ram_c_21_0_enable)
  );

  wire [20-1:0] ram_c_22_0_addr;
  wire [32-1:0] ram_c_22_0_rdata;
  wire [32-1:0] ram_c_22_0_wdata;
  wire ram_c_22_0_wenable;
  wire ram_c_22_0_enable;

  ram_c_22
  inst_ram_c_22
  (
    .CLK(CLK),
    .ram_c_22_0_addr(ram_c_22_0_addr),
    .ram_c_22_0_rdata(ram_c_22_0_rdata),
    .ram_c_22_0_wdata(ram_c_22_0_wdata),
    .ram_c_22_0_wenable(ram_c_22_0_wenable),
    .ram_c_22_0_enable(ram_c_22_0_enable)
  );

  wire [20-1:0] ram_c_23_0_addr;
  wire [32-1:0] ram_c_23_0_rdata;
  wire [32-1:0] ram_c_23_0_wdata;
  wire ram_c_23_0_wenable;
  wire ram_c_23_0_enable;

  ram_c_23
  inst_ram_c_23
  (
    .CLK(CLK),
    .ram_c_23_0_addr(ram_c_23_0_addr),
    .ram_c_23_0_rdata(ram_c_23_0_rdata),
    .ram_c_23_0_wdata(ram_c_23_0_wdata),
    .ram_c_23_0_wenable(ram_c_23_0_wenable),
    .ram_c_23_0_enable(ram_c_23_0_enable)
  );

  wire [20-1:0] ram_c_24_0_addr;
  wire [32-1:0] ram_c_24_0_rdata;
  wire [32-1:0] ram_c_24_0_wdata;
  wire ram_c_24_0_wenable;
  wire ram_c_24_0_enable;

  ram_c_24
  inst_ram_c_24
  (
    .CLK(CLK),
    .ram_c_24_0_addr(ram_c_24_0_addr),
    .ram_c_24_0_rdata(ram_c_24_0_rdata),
    .ram_c_24_0_wdata(ram_c_24_0_wdata),
    .ram_c_24_0_wenable(ram_c_24_0_wenable),
    .ram_c_24_0_enable(ram_c_24_0_enable)
  );

  wire [20-1:0] ram_c_25_0_addr;
  wire [32-1:0] ram_c_25_0_rdata;
  wire [32-1:0] ram_c_25_0_wdata;
  wire ram_c_25_0_wenable;
  wire ram_c_25_0_enable;

  ram_c_25
  inst_ram_c_25
  (
    .CLK(CLK),
    .ram_c_25_0_addr(ram_c_25_0_addr),
    .ram_c_25_0_rdata(ram_c_25_0_rdata),
    .ram_c_25_0_wdata(ram_c_25_0_wdata),
    .ram_c_25_0_wenable(ram_c_25_0_wenable),
    .ram_c_25_0_enable(ram_c_25_0_enable)
  );

  wire [20-1:0] ram_c_26_0_addr;
  wire [32-1:0] ram_c_26_0_rdata;
  wire [32-1:0] ram_c_26_0_wdata;
  wire ram_c_26_0_wenable;
  wire ram_c_26_0_enable;

  ram_c_26
  inst_ram_c_26
  (
    .CLK(CLK),
    .ram_c_26_0_addr(ram_c_26_0_addr),
    .ram_c_26_0_rdata(ram_c_26_0_rdata),
    .ram_c_26_0_wdata(ram_c_26_0_wdata),
    .ram_c_26_0_wenable(ram_c_26_0_wenable),
    .ram_c_26_0_enable(ram_c_26_0_enable)
  );

  wire [20-1:0] ram_c_27_0_addr;
  wire [32-1:0] ram_c_27_0_rdata;
  wire [32-1:0] ram_c_27_0_wdata;
  wire ram_c_27_0_wenable;
  wire ram_c_27_0_enable;

  ram_c_27
  inst_ram_c_27
  (
    .CLK(CLK),
    .ram_c_27_0_addr(ram_c_27_0_addr),
    .ram_c_27_0_rdata(ram_c_27_0_rdata),
    .ram_c_27_0_wdata(ram_c_27_0_wdata),
    .ram_c_27_0_wenable(ram_c_27_0_wenable),
    .ram_c_27_0_enable(ram_c_27_0_enable)
  );

  wire [20-1:0] ram_c_28_0_addr;
  wire [32-1:0] ram_c_28_0_rdata;
  wire [32-1:0] ram_c_28_0_wdata;
  wire ram_c_28_0_wenable;
  wire ram_c_28_0_enable;

  ram_c_28
  inst_ram_c_28
  (
    .CLK(CLK),
    .ram_c_28_0_addr(ram_c_28_0_addr),
    .ram_c_28_0_rdata(ram_c_28_0_rdata),
    .ram_c_28_0_wdata(ram_c_28_0_wdata),
    .ram_c_28_0_wenable(ram_c_28_0_wenable),
    .ram_c_28_0_enable(ram_c_28_0_enable)
  );

  wire [20-1:0] ram_c_29_0_addr;
  wire [32-1:0] ram_c_29_0_rdata;
  wire [32-1:0] ram_c_29_0_wdata;
  wire ram_c_29_0_wenable;
  wire ram_c_29_0_enable;

  ram_c_29
  inst_ram_c_29
  (
    .CLK(CLK),
    .ram_c_29_0_addr(ram_c_29_0_addr),
    .ram_c_29_0_rdata(ram_c_29_0_rdata),
    .ram_c_29_0_wdata(ram_c_29_0_wdata),
    .ram_c_29_0_wenable(ram_c_29_0_wenable),
    .ram_c_29_0_enable(ram_c_29_0_enable)
  );

  wire [20-1:0] ram_c_30_0_addr;
  wire [32-1:0] ram_c_30_0_rdata;
  wire [32-1:0] ram_c_30_0_wdata;
  wire ram_c_30_0_wenable;
  wire ram_c_30_0_enable;

  ram_c_30
  inst_ram_c_30
  (
    .CLK(CLK),
    .ram_c_30_0_addr(ram_c_30_0_addr),
    .ram_c_30_0_rdata(ram_c_30_0_rdata),
    .ram_c_30_0_wdata(ram_c_30_0_wdata),
    .ram_c_30_0_wenable(ram_c_30_0_wenable),
    .ram_c_30_0_enable(ram_c_30_0_enable)
  );

  wire [20-1:0] ram_c_31_0_addr;
  wire [32-1:0] ram_c_31_0_rdata;
  wire [32-1:0] ram_c_31_0_wdata;
  wire ram_c_31_0_wenable;
  wire ram_c_31_0_enable;

  ram_c_31
  inst_ram_c_31
  (
    .CLK(CLK),
    .ram_c_31_0_addr(ram_c_31_0_addr),
    .ram_c_31_0_rdata(ram_c_31_0_rdata),
    .ram_c_31_0_wdata(ram_c_31_0_wdata),
    .ram_c_31_0_wenable(ram_c_31_0_wenable),
    .ram_c_31_0_enable(ram_c_31_0_enable)
  );

  wire [20-1:0] ram_x_0_addr;
  wire [32-1:0] ram_x_0_rdata;
  wire [32-1:0] ram_x_0_wdata;
  wire ram_x_0_wenable;
  wire ram_x_0_enable;

  ram_x
  inst_ram_x
  (
    .CLK(CLK),
    .ram_x_0_addr(ram_x_0_addr),
    .ram_x_0_rdata(ram_x_0_rdata),
    .ram_x_0_wdata(ram_x_0_wdata),
    .ram_x_0_wenable(ram_x_0_wenable),
    .ram_x_0_enable(ram_x_0_enable)
  );

  wire [20-1:0] ram_y_0_addr;
  wire [32-1:0] ram_y_0_rdata;
  wire [32-1:0] ram_y_0_wdata;
  wire ram_y_0_wenable;
  wire ram_y_0_enable;

  ram_y
  inst_ram_y
  (
    .CLK(CLK),
    .ram_y_0_addr(ram_y_0_addr),
    .ram_y_0_rdata(ram_y_0_rdata),
    .ram_y_0_wdata(ram_y_0_wdata),
    .ram_y_0_wenable(ram_y_0_wenable),
    .ram_y_0_enable(ram_y_0_enable)
  );

  wire [20-1:0] ram_z_0_addr;
  wire [32-1:0] ram_z_0_rdata;
  wire [32-1:0] ram_z_0_wdata;
  wire ram_z_0_wenable;
  wire ram_z_0_enable;

  ram_z
  inst_ram_z
  (
    .CLK(CLK),
    .ram_z_0_addr(ram_z_0_addr),
    .ram_z_0_rdata(ram_z_0_rdata),
    .ram_z_0_wdata(ram_z_0_wdata),
    .ram_z_0_wenable(ram_z_0_wenable),
    .ram_z_0_enable(ram_z_0_enable)
  );

  reg _mystream_stream_ivalid;
  wire _mystream_stream_oready;
  wire _mystream_stream_internal_oready;
  assign _mystream_stream_internal_oready = 1;
  assign _mystream_stream_oready = _mystream_stream_internal_oready;
  reg [32-1:0] _mystream_fsm;
  localparam _mystream_fsm_init = 0;
  wire _mystream_run_flag;
  reg _mystream_source_start;
  wire _mystream_source_stop;
  reg _mystream_source_busy;
  wire _mystream_sink_start;
  wire _mystream_sink_stop;
  wire _mystream_sink_busy;
  wire _mystream_busy;
  reg _mystream_busy_reg;
  wire _mystream_is_root;
  assign _mystream_is_root = 1;
  reg [32-1:0] _mystream_size_next_parameter_data;
  reg [32-1:0] _mystream_tensor_size_next_parameter_data;
  reg _mystream_a0_idle;
  reg [33-1:0] _mystream_a0_source_count;
  reg [5-1:0] _mystream_a0_source_mode;
  reg [16-1:0] _mystream_a0_source_generator_id;
  reg [32-1:0] _mystream_a0_source_offset;
  reg [33-1:0] _mystream_a0_source_size;
  reg [32-1:0] _mystream_a0_source_stride;
  reg [32-1:0] _mystream_a0_source_offset_buf;
  reg [33-1:0] _mystream_a0_source_size_buf;
  reg [32-1:0] _mystream_a0_source_stride_buf;
  reg [8-1:0] _mystream_a0_source_sel;
  reg [32-1:0] _mystream_a0_source_ram_raddr;
  reg _mystream_a0_source_ram_renable;
  wire [32-1:0] _mystream_a0_source_ram_rdata;
  reg _mystream_a0_source_fifo_deq;
  wire [32-1:0] _mystream_a0_source_fifo_rdata;
  reg [32-1:0] _mystream_a0_source_empty_data;
  reg _mystream_a1_idle;
  reg [33-1:0] _mystream_a1_source_count;
  reg [5-1:0] _mystream_a1_source_mode;
  reg [16-1:0] _mystream_a1_source_generator_id;
  reg [32-1:0] _mystream_a1_source_offset;
  reg [33-1:0] _mystream_a1_source_size;
  reg [32-1:0] _mystream_a1_source_stride;
  reg [32-1:0] _mystream_a1_source_offset_buf;
  reg [33-1:0] _mystream_a1_source_size_buf;
  reg [32-1:0] _mystream_a1_source_stride_buf;
  reg [8-1:0] _mystream_a1_source_sel;
  reg [32-1:0] _mystream_a1_source_ram_raddr;
  reg _mystream_a1_source_ram_renable;
  wire [32-1:0] _mystream_a1_source_ram_rdata;
  reg _mystream_a1_source_fifo_deq;
  wire [32-1:0] _mystream_a1_source_fifo_rdata;
  reg [32-1:0] _mystream_a1_source_empty_data;
  reg _mystream_a2_idle;
  reg [33-1:0] _mystream_a2_source_count;
  reg [5-1:0] _mystream_a2_source_mode;
  reg [16-1:0] _mystream_a2_source_generator_id;
  reg [32-1:0] _mystream_a2_source_offset;
  reg [33-1:0] _mystream_a2_source_size;
  reg [32-1:0] _mystream_a2_source_stride;
  reg [32-1:0] _mystream_a2_source_offset_buf;
  reg [33-1:0] _mystream_a2_source_size_buf;
  reg [32-1:0] _mystream_a2_source_stride_buf;
  reg [8-1:0] _mystream_a2_source_sel;
  reg [32-1:0] _mystream_a2_source_ram_raddr;
  reg _mystream_a2_source_ram_renable;
  wire [32-1:0] _mystream_a2_source_ram_rdata;
  reg _mystream_a2_source_fifo_deq;
  wire [32-1:0] _mystream_a2_source_fifo_rdata;
  reg [32-1:0] _mystream_a2_source_empty_data;
  reg _mystream_a3_idle;
  reg [33-1:0] _mystream_a3_source_count;
  reg [5-1:0] _mystream_a3_source_mode;
  reg [16-1:0] _mystream_a3_source_generator_id;
  reg [32-1:0] _mystream_a3_source_offset;
  reg [33-1:0] _mystream_a3_source_size;
  reg [32-1:0] _mystream_a3_source_stride;
  reg [32-1:0] _mystream_a3_source_offset_buf;
  reg [33-1:0] _mystream_a3_source_size_buf;
  reg [32-1:0] _mystream_a3_source_stride_buf;
  reg [8-1:0] _mystream_a3_source_sel;
  reg [32-1:0] _mystream_a3_source_ram_raddr;
  reg _mystream_a3_source_ram_renable;
  wire [32-1:0] _mystream_a3_source_ram_rdata;
  reg _mystream_a3_source_fifo_deq;
  wire [32-1:0] _mystream_a3_source_fifo_rdata;
  reg [32-1:0] _mystream_a3_source_empty_data;
  reg _mystream_a4_idle;
  reg [33-1:0] _mystream_a4_source_count;
  reg [5-1:0] _mystream_a4_source_mode;
  reg [16-1:0] _mystream_a4_source_generator_id;
  reg [32-1:0] _mystream_a4_source_offset;
  reg [33-1:0] _mystream_a4_source_size;
  reg [32-1:0] _mystream_a4_source_stride;
  reg [32-1:0] _mystream_a4_source_offset_buf;
  reg [33-1:0] _mystream_a4_source_size_buf;
  reg [32-1:0] _mystream_a4_source_stride_buf;
  reg [8-1:0] _mystream_a4_source_sel;
  reg [32-1:0] _mystream_a4_source_ram_raddr;
  reg _mystream_a4_source_ram_renable;
  wire [32-1:0] _mystream_a4_source_ram_rdata;
  reg _mystream_a4_source_fifo_deq;
  wire [32-1:0] _mystream_a4_source_fifo_rdata;
  reg [32-1:0] _mystream_a4_source_empty_data;
  reg _mystream_a5_idle;
  reg [33-1:0] _mystream_a5_source_count;
  reg [5-1:0] _mystream_a5_source_mode;
  reg [16-1:0] _mystream_a5_source_generator_id;
  reg [32-1:0] _mystream_a5_source_offset;
  reg [33-1:0] _mystream_a5_source_size;
  reg [32-1:0] _mystream_a5_source_stride;
  reg [32-1:0] _mystream_a5_source_offset_buf;
  reg [33-1:0] _mystream_a5_source_size_buf;
  reg [32-1:0] _mystream_a5_source_stride_buf;
  reg [8-1:0] _mystream_a5_source_sel;
  reg [32-1:0] _mystream_a5_source_ram_raddr;
  reg _mystream_a5_source_ram_renable;
  wire [32-1:0] _mystream_a5_source_ram_rdata;
  reg _mystream_a5_source_fifo_deq;
  wire [32-1:0] _mystream_a5_source_fifo_rdata;
  reg [32-1:0] _mystream_a5_source_empty_data;
  reg _mystream_a6_idle;
  reg [33-1:0] _mystream_a6_source_count;
  reg [5-1:0] _mystream_a6_source_mode;
  reg [16-1:0] _mystream_a6_source_generator_id;
  reg [32-1:0] _mystream_a6_source_offset;
  reg [33-1:0] _mystream_a6_source_size;
  reg [32-1:0] _mystream_a6_source_stride;
  reg [32-1:0] _mystream_a6_source_offset_buf;
  reg [33-1:0] _mystream_a6_source_size_buf;
  reg [32-1:0] _mystream_a6_source_stride_buf;
  reg [8-1:0] _mystream_a6_source_sel;
  reg [32-1:0] _mystream_a6_source_ram_raddr;
  reg _mystream_a6_source_ram_renable;
  wire [32-1:0] _mystream_a6_source_ram_rdata;
  reg _mystream_a6_source_fifo_deq;
  wire [32-1:0] _mystream_a6_source_fifo_rdata;
  reg [32-1:0] _mystream_a6_source_empty_data;
  reg _mystream_a7_idle;
  reg [33-1:0] _mystream_a7_source_count;
  reg [5-1:0] _mystream_a7_source_mode;
  reg [16-1:0] _mystream_a7_source_generator_id;
  reg [32-1:0] _mystream_a7_source_offset;
  reg [33-1:0] _mystream_a7_source_size;
  reg [32-1:0] _mystream_a7_source_stride;
  reg [32-1:0] _mystream_a7_source_offset_buf;
  reg [33-1:0] _mystream_a7_source_size_buf;
  reg [32-1:0] _mystream_a7_source_stride_buf;
  reg [8-1:0] _mystream_a7_source_sel;
  reg [32-1:0] _mystream_a7_source_ram_raddr;
  reg _mystream_a7_source_ram_renable;
  wire [32-1:0] _mystream_a7_source_ram_rdata;
  reg _mystream_a7_source_fifo_deq;
  wire [32-1:0] _mystream_a7_source_fifo_rdata;
  reg [32-1:0] _mystream_a7_source_empty_data;
  reg _mystream_a8_idle;
  reg [33-1:0] _mystream_a8_source_count;
  reg [5-1:0] _mystream_a8_source_mode;
  reg [16-1:0] _mystream_a8_source_generator_id;
  reg [32-1:0] _mystream_a8_source_offset;
  reg [33-1:0] _mystream_a8_source_size;
  reg [32-1:0] _mystream_a8_source_stride;
  reg [32-1:0] _mystream_a8_source_offset_buf;
  reg [33-1:0] _mystream_a8_source_size_buf;
  reg [32-1:0] _mystream_a8_source_stride_buf;
  reg [8-1:0] _mystream_a8_source_sel;
  reg [32-1:0] _mystream_a8_source_ram_raddr;
  reg _mystream_a8_source_ram_renable;
  wire [32-1:0] _mystream_a8_source_ram_rdata;
  reg _mystream_a8_source_fifo_deq;
  wire [32-1:0] _mystream_a8_source_fifo_rdata;
  reg [32-1:0] _mystream_a8_source_empty_data;
  reg _mystream_a9_idle;
  reg [33-1:0] _mystream_a9_source_count;
  reg [5-1:0] _mystream_a9_source_mode;
  reg [16-1:0] _mystream_a9_source_generator_id;
  reg [32-1:0] _mystream_a9_source_offset;
  reg [33-1:0] _mystream_a9_source_size;
  reg [32-1:0] _mystream_a9_source_stride;
  reg [32-1:0] _mystream_a9_source_offset_buf;
  reg [33-1:0] _mystream_a9_source_size_buf;
  reg [32-1:0] _mystream_a9_source_stride_buf;
  reg [8-1:0] _mystream_a9_source_sel;
  reg [32-1:0] _mystream_a9_source_ram_raddr;
  reg _mystream_a9_source_ram_renable;
  wire [32-1:0] _mystream_a9_source_ram_rdata;
  reg _mystream_a9_source_fifo_deq;
  wire [32-1:0] _mystream_a9_source_fifo_rdata;
  reg [32-1:0] _mystream_a9_source_empty_data;
  reg _mystream_a10_idle;
  reg [33-1:0] _mystream_a10_source_count;
  reg [5-1:0] _mystream_a10_source_mode;
  reg [16-1:0] _mystream_a10_source_generator_id;
  reg [32-1:0] _mystream_a10_source_offset;
  reg [33-1:0] _mystream_a10_source_size;
  reg [32-1:0] _mystream_a10_source_stride;
  reg [32-1:0] _mystream_a10_source_offset_buf;
  reg [33-1:0] _mystream_a10_source_size_buf;
  reg [32-1:0] _mystream_a10_source_stride_buf;
  reg [8-1:0] _mystream_a10_source_sel;
  reg [32-1:0] _mystream_a10_source_ram_raddr;
  reg _mystream_a10_source_ram_renable;
  wire [32-1:0] _mystream_a10_source_ram_rdata;
  reg _mystream_a10_source_fifo_deq;
  wire [32-1:0] _mystream_a10_source_fifo_rdata;
  reg [32-1:0] _mystream_a10_source_empty_data;
  reg _mystream_a11_idle;
  reg [33-1:0] _mystream_a11_source_count;
  reg [5-1:0] _mystream_a11_source_mode;
  reg [16-1:0] _mystream_a11_source_generator_id;
  reg [32-1:0] _mystream_a11_source_offset;
  reg [33-1:0] _mystream_a11_source_size;
  reg [32-1:0] _mystream_a11_source_stride;
  reg [32-1:0] _mystream_a11_source_offset_buf;
  reg [33-1:0] _mystream_a11_source_size_buf;
  reg [32-1:0] _mystream_a11_source_stride_buf;
  reg [8-1:0] _mystream_a11_source_sel;
  reg [32-1:0] _mystream_a11_source_ram_raddr;
  reg _mystream_a11_source_ram_renable;
  wire [32-1:0] _mystream_a11_source_ram_rdata;
  reg _mystream_a11_source_fifo_deq;
  wire [32-1:0] _mystream_a11_source_fifo_rdata;
  reg [32-1:0] _mystream_a11_source_empty_data;
  reg _mystream_a12_idle;
  reg [33-1:0] _mystream_a12_source_count;
  reg [5-1:0] _mystream_a12_source_mode;
  reg [16-1:0] _mystream_a12_source_generator_id;
  reg [32-1:0] _mystream_a12_source_offset;
  reg [33-1:0] _mystream_a12_source_size;
  reg [32-1:0] _mystream_a12_source_stride;
  reg [32-1:0] _mystream_a12_source_offset_buf;
  reg [33-1:0] _mystream_a12_source_size_buf;
  reg [32-1:0] _mystream_a12_source_stride_buf;
  reg [8-1:0] _mystream_a12_source_sel;
  reg [32-1:0] _mystream_a12_source_ram_raddr;
  reg _mystream_a12_source_ram_renable;
  wire [32-1:0] _mystream_a12_source_ram_rdata;
  reg _mystream_a12_source_fifo_deq;
  wire [32-1:0] _mystream_a12_source_fifo_rdata;
  reg [32-1:0] _mystream_a12_source_empty_data;
  reg _mystream_a13_idle;
  reg [33-1:0] _mystream_a13_source_count;
  reg [5-1:0] _mystream_a13_source_mode;
  reg [16-1:0] _mystream_a13_source_generator_id;
  reg [32-1:0] _mystream_a13_source_offset;
  reg [33-1:0] _mystream_a13_source_size;
  reg [32-1:0] _mystream_a13_source_stride;
  reg [32-1:0] _mystream_a13_source_offset_buf;
  reg [33-1:0] _mystream_a13_source_size_buf;
  reg [32-1:0] _mystream_a13_source_stride_buf;
  reg [8-1:0] _mystream_a13_source_sel;
  reg [32-1:0] _mystream_a13_source_ram_raddr;
  reg _mystream_a13_source_ram_renable;
  wire [32-1:0] _mystream_a13_source_ram_rdata;
  reg _mystream_a13_source_fifo_deq;
  wire [32-1:0] _mystream_a13_source_fifo_rdata;
  reg [32-1:0] _mystream_a13_source_empty_data;
  reg _mystream_a14_idle;
  reg [33-1:0] _mystream_a14_source_count;
  reg [5-1:0] _mystream_a14_source_mode;
  reg [16-1:0] _mystream_a14_source_generator_id;
  reg [32-1:0] _mystream_a14_source_offset;
  reg [33-1:0] _mystream_a14_source_size;
  reg [32-1:0] _mystream_a14_source_stride;
  reg [32-1:0] _mystream_a14_source_offset_buf;
  reg [33-1:0] _mystream_a14_source_size_buf;
  reg [32-1:0] _mystream_a14_source_stride_buf;
  reg [8-1:0] _mystream_a14_source_sel;
  reg [32-1:0] _mystream_a14_source_ram_raddr;
  reg _mystream_a14_source_ram_renable;
  wire [32-1:0] _mystream_a14_source_ram_rdata;
  reg _mystream_a14_source_fifo_deq;
  wire [32-1:0] _mystream_a14_source_fifo_rdata;
  reg [32-1:0] _mystream_a14_source_empty_data;
  reg _mystream_a15_idle;
  reg [33-1:0] _mystream_a15_source_count;
  reg [5-1:0] _mystream_a15_source_mode;
  reg [16-1:0] _mystream_a15_source_generator_id;
  reg [32-1:0] _mystream_a15_source_offset;
  reg [33-1:0] _mystream_a15_source_size;
  reg [32-1:0] _mystream_a15_source_stride;
  reg [32-1:0] _mystream_a15_source_offset_buf;
  reg [33-1:0] _mystream_a15_source_size_buf;
  reg [32-1:0] _mystream_a15_source_stride_buf;
  reg [8-1:0] _mystream_a15_source_sel;
  reg [32-1:0] _mystream_a15_source_ram_raddr;
  reg _mystream_a15_source_ram_renable;
  wire [32-1:0] _mystream_a15_source_ram_rdata;
  reg _mystream_a15_source_fifo_deq;
  wire [32-1:0] _mystream_a15_source_fifo_rdata;
  reg [32-1:0] _mystream_a15_source_empty_data;
  reg _mystream_a16_idle;
  reg [33-1:0] _mystream_a16_source_count;
  reg [5-1:0] _mystream_a16_source_mode;
  reg [16-1:0] _mystream_a16_source_generator_id;
  reg [32-1:0] _mystream_a16_source_offset;
  reg [33-1:0] _mystream_a16_source_size;
  reg [32-1:0] _mystream_a16_source_stride;
  reg [32-1:0] _mystream_a16_source_offset_buf;
  reg [33-1:0] _mystream_a16_source_size_buf;
  reg [32-1:0] _mystream_a16_source_stride_buf;
  reg [8-1:0] _mystream_a16_source_sel;
  reg [32-1:0] _mystream_a16_source_ram_raddr;
  reg _mystream_a16_source_ram_renable;
  wire [32-1:0] _mystream_a16_source_ram_rdata;
  reg _mystream_a16_source_fifo_deq;
  wire [32-1:0] _mystream_a16_source_fifo_rdata;
  reg [32-1:0] _mystream_a16_source_empty_data;
  reg _mystream_a17_idle;
  reg [33-1:0] _mystream_a17_source_count;
  reg [5-1:0] _mystream_a17_source_mode;
  reg [16-1:0] _mystream_a17_source_generator_id;
  reg [32-1:0] _mystream_a17_source_offset;
  reg [33-1:0] _mystream_a17_source_size;
  reg [32-1:0] _mystream_a17_source_stride;
  reg [32-1:0] _mystream_a17_source_offset_buf;
  reg [33-1:0] _mystream_a17_source_size_buf;
  reg [32-1:0] _mystream_a17_source_stride_buf;
  reg [8-1:0] _mystream_a17_source_sel;
  reg [32-1:0] _mystream_a17_source_ram_raddr;
  reg _mystream_a17_source_ram_renable;
  wire [32-1:0] _mystream_a17_source_ram_rdata;
  reg _mystream_a17_source_fifo_deq;
  wire [32-1:0] _mystream_a17_source_fifo_rdata;
  reg [32-1:0] _mystream_a17_source_empty_data;
  reg _mystream_a18_idle;
  reg [33-1:0] _mystream_a18_source_count;
  reg [5-1:0] _mystream_a18_source_mode;
  reg [16-1:0] _mystream_a18_source_generator_id;
  reg [32-1:0] _mystream_a18_source_offset;
  reg [33-1:0] _mystream_a18_source_size;
  reg [32-1:0] _mystream_a18_source_stride;
  reg [32-1:0] _mystream_a18_source_offset_buf;
  reg [33-1:0] _mystream_a18_source_size_buf;
  reg [32-1:0] _mystream_a18_source_stride_buf;
  reg [8-1:0] _mystream_a18_source_sel;
  reg [32-1:0] _mystream_a18_source_ram_raddr;
  reg _mystream_a18_source_ram_renable;
  wire [32-1:0] _mystream_a18_source_ram_rdata;
  reg _mystream_a18_source_fifo_deq;
  wire [32-1:0] _mystream_a18_source_fifo_rdata;
  reg [32-1:0] _mystream_a18_source_empty_data;
  reg _mystream_a19_idle;
  reg [33-1:0] _mystream_a19_source_count;
  reg [5-1:0] _mystream_a19_source_mode;
  reg [16-1:0] _mystream_a19_source_generator_id;
  reg [32-1:0] _mystream_a19_source_offset;
  reg [33-1:0] _mystream_a19_source_size;
  reg [32-1:0] _mystream_a19_source_stride;
  reg [32-1:0] _mystream_a19_source_offset_buf;
  reg [33-1:0] _mystream_a19_source_size_buf;
  reg [32-1:0] _mystream_a19_source_stride_buf;
  reg [8-1:0] _mystream_a19_source_sel;
  reg [32-1:0] _mystream_a19_source_ram_raddr;
  reg _mystream_a19_source_ram_renable;
  wire [32-1:0] _mystream_a19_source_ram_rdata;
  reg _mystream_a19_source_fifo_deq;
  wire [32-1:0] _mystream_a19_source_fifo_rdata;
  reg [32-1:0] _mystream_a19_source_empty_data;
  reg _mystream_a20_idle;
  reg [33-1:0] _mystream_a20_source_count;
  reg [5-1:0] _mystream_a20_source_mode;
  reg [16-1:0] _mystream_a20_source_generator_id;
  reg [32-1:0] _mystream_a20_source_offset;
  reg [33-1:0] _mystream_a20_source_size;
  reg [32-1:0] _mystream_a20_source_stride;
  reg [32-1:0] _mystream_a20_source_offset_buf;
  reg [33-1:0] _mystream_a20_source_size_buf;
  reg [32-1:0] _mystream_a20_source_stride_buf;
  reg [8-1:0] _mystream_a20_source_sel;
  reg [32-1:0] _mystream_a20_source_ram_raddr;
  reg _mystream_a20_source_ram_renable;
  wire [32-1:0] _mystream_a20_source_ram_rdata;
  reg _mystream_a20_source_fifo_deq;
  wire [32-1:0] _mystream_a20_source_fifo_rdata;
  reg [32-1:0] _mystream_a20_source_empty_data;
  reg _mystream_a21_idle;
  reg [33-1:0] _mystream_a21_source_count;
  reg [5-1:0] _mystream_a21_source_mode;
  reg [16-1:0] _mystream_a21_source_generator_id;
  reg [32-1:0] _mystream_a21_source_offset;
  reg [33-1:0] _mystream_a21_source_size;
  reg [32-1:0] _mystream_a21_source_stride;
  reg [32-1:0] _mystream_a21_source_offset_buf;
  reg [33-1:0] _mystream_a21_source_size_buf;
  reg [32-1:0] _mystream_a21_source_stride_buf;
  reg [8-1:0] _mystream_a21_source_sel;
  reg [32-1:0] _mystream_a21_source_ram_raddr;
  reg _mystream_a21_source_ram_renable;
  wire [32-1:0] _mystream_a21_source_ram_rdata;
  reg _mystream_a21_source_fifo_deq;
  wire [32-1:0] _mystream_a21_source_fifo_rdata;
  reg [32-1:0] _mystream_a21_source_empty_data;
  reg _mystream_a22_idle;
  reg [33-1:0] _mystream_a22_source_count;
  reg [5-1:0] _mystream_a22_source_mode;
  reg [16-1:0] _mystream_a22_source_generator_id;
  reg [32-1:0] _mystream_a22_source_offset;
  reg [33-1:0] _mystream_a22_source_size;
  reg [32-1:0] _mystream_a22_source_stride;
  reg [32-1:0] _mystream_a22_source_offset_buf;
  reg [33-1:0] _mystream_a22_source_size_buf;
  reg [32-1:0] _mystream_a22_source_stride_buf;
  reg [8-1:0] _mystream_a22_source_sel;
  reg [32-1:0] _mystream_a22_source_ram_raddr;
  reg _mystream_a22_source_ram_renable;
  wire [32-1:0] _mystream_a22_source_ram_rdata;
  reg _mystream_a22_source_fifo_deq;
  wire [32-1:0] _mystream_a22_source_fifo_rdata;
  reg [32-1:0] _mystream_a22_source_empty_data;
  reg _mystream_a23_idle;
  reg [33-1:0] _mystream_a23_source_count;
  reg [5-1:0] _mystream_a23_source_mode;
  reg [16-1:0] _mystream_a23_source_generator_id;
  reg [32-1:0] _mystream_a23_source_offset;
  reg [33-1:0] _mystream_a23_source_size;
  reg [32-1:0] _mystream_a23_source_stride;
  reg [32-1:0] _mystream_a23_source_offset_buf;
  reg [33-1:0] _mystream_a23_source_size_buf;
  reg [32-1:0] _mystream_a23_source_stride_buf;
  reg [8-1:0] _mystream_a23_source_sel;
  reg [32-1:0] _mystream_a23_source_ram_raddr;
  reg _mystream_a23_source_ram_renable;
  wire [32-1:0] _mystream_a23_source_ram_rdata;
  reg _mystream_a23_source_fifo_deq;
  wire [32-1:0] _mystream_a23_source_fifo_rdata;
  reg [32-1:0] _mystream_a23_source_empty_data;
  reg _mystream_a24_idle;
  reg [33-1:0] _mystream_a24_source_count;
  reg [5-1:0] _mystream_a24_source_mode;
  reg [16-1:0] _mystream_a24_source_generator_id;
  reg [32-1:0] _mystream_a24_source_offset;
  reg [33-1:0] _mystream_a24_source_size;
  reg [32-1:0] _mystream_a24_source_stride;
  reg [32-1:0] _mystream_a24_source_offset_buf;
  reg [33-1:0] _mystream_a24_source_size_buf;
  reg [32-1:0] _mystream_a24_source_stride_buf;
  reg [8-1:0] _mystream_a24_source_sel;
  reg [32-1:0] _mystream_a24_source_ram_raddr;
  reg _mystream_a24_source_ram_renable;
  wire [32-1:0] _mystream_a24_source_ram_rdata;
  reg _mystream_a24_source_fifo_deq;
  wire [32-1:0] _mystream_a24_source_fifo_rdata;
  reg [32-1:0] _mystream_a24_source_empty_data;
  reg _mystream_a25_idle;
  reg [33-1:0] _mystream_a25_source_count;
  reg [5-1:0] _mystream_a25_source_mode;
  reg [16-1:0] _mystream_a25_source_generator_id;
  reg [32-1:0] _mystream_a25_source_offset;
  reg [33-1:0] _mystream_a25_source_size;
  reg [32-1:0] _mystream_a25_source_stride;
  reg [32-1:0] _mystream_a25_source_offset_buf;
  reg [33-1:0] _mystream_a25_source_size_buf;
  reg [32-1:0] _mystream_a25_source_stride_buf;
  reg [8-1:0] _mystream_a25_source_sel;
  reg [32-1:0] _mystream_a25_source_ram_raddr;
  reg _mystream_a25_source_ram_renable;
  wire [32-1:0] _mystream_a25_source_ram_rdata;
  reg _mystream_a25_source_fifo_deq;
  wire [32-1:0] _mystream_a25_source_fifo_rdata;
  reg [32-1:0] _mystream_a25_source_empty_data;
  reg _mystream_a26_idle;
  reg [33-1:0] _mystream_a26_source_count;
  reg [5-1:0] _mystream_a26_source_mode;
  reg [16-1:0] _mystream_a26_source_generator_id;
  reg [32-1:0] _mystream_a26_source_offset;
  reg [33-1:0] _mystream_a26_source_size;
  reg [32-1:0] _mystream_a26_source_stride;
  reg [32-1:0] _mystream_a26_source_offset_buf;
  reg [33-1:0] _mystream_a26_source_size_buf;
  reg [32-1:0] _mystream_a26_source_stride_buf;
  reg [8-1:0] _mystream_a26_source_sel;
  reg [32-1:0] _mystream_a26_source_ram_raddr;
  reg _mystream_a26_source_ram_renable;
  wire [32-1:0] _mystream_a26_source_ram_rdata;
  reg _mystream_a26_source_fifo_deq;
  wire [32-1:0] _mystream_a26_source_fifo_rdata;
  reg [32-1:0] _mystream_a26_source_empty_data;
  reg _mystream_a27_idle;
  reg [33-1:0] _mystream_a27_source_count;
  reg [5-1:0] _mystream_a27_source_mode;
  reg [16-1:0] _mystream_a27_source_generator_id;
  reg [32-1:0] _mystream_a27_source_offset;
  reg [33-1:0] _mystream_a27_source_size;
  reg [32-1:0] _mystream_a27_source_stride;
  reg [32-1:0] _mystream_a27_source_offset_buf;
  reg [33-1:0] _mystream_a27_source_size_buf;
  reg [32-1:0] _mystream_a27_source_stride_buf;
  reg [8-1:0] _mystream_a27_source_sel;
  reg [32-1:0] _mystream_a27_source_ram_raddr;
  reg _mystream_a27_source_ram_renable;
  wire [32-1:0] _mystream_a27_source_ram_rdata;
  reg _mystream_a27_source_fifo_deq;
  wire [32-1:0] _mystream_a27_source_fifo_rdata;
  reg [32-1:0] _mystream_a27_source_empty_data;
  reg _mystream_a28_idle;
  reg [33-1:0] _mystream_a28_source_count;
  reg [5-1:0] _mystream_a28_source_mode;
  reg [16-1:0] _mystream_a28_source_generator_id;
  reg [32-1:0] _mystream_a28_source_offset;
  reg [33-1:0] _mystream_a28_source_size;
  reg [32-1:0] _mystream_a28_source_stride;
  reg [32-1:0] _mystream_a28_source_offset_buf;
  reg [33-1:0] _mystream_a28_source_size_buf;
  reg [32-1:0] _mystream_a28_source_stride_buf;
  reg [8-1:0] _mystream_a28_source_sel;
  reg [32-1:0] _mystream_a28_source_ram_raddr;
  reg _mystream_a28_source_ram_renable;
  wire [32-1:0] _mystream_a28_source_ram_rdata;
  reg _mystream_a28_source_fifo_deq;
  wire [32-1:0] _mystream_a28_source_fifo_rdata;
  reg [32-1:0] _mystream_a28_source_empty_data;
  reg _mystream_a29_idle;
  reg [33-1:0] _mystream_a29_source_count;
  reg [5-1:0] _mystream_a29_source_mode;
  reg [16-1:0] _mystream_a29_source_generator_id;
  reg [32-1:0] _mystream_a29_source_offset;
  reg [33-1:0] _mystream_a29_source_size;
  reg [32-1:0] _mystream_a29_source_stride;
  reg [32-1:0] _mystream_a29_source_offset_buf;
  reg [33-1:0] _mystream_a29_source_size_buf;
  reg [32-1:0] _mystream_a29_source_stride_buf;
  reg [8-1:0] _mystream_a29_source_sel;
  reg [32-1:0] _mystream_a29_source_ram_raddr;
  reg _mystream_a29_source_ram_renable;
  wire [32-1:0] _mystream_a29_source_ram_rdata;
  reg _mystream_a29_source_fifo_deq;
  wire [32-1:0] _mystream_a29_source_fifo_rdata;
  reg [32-1:0] _mystream_a29_source_empty_data;
  reg _mystream_a30_idle;
  reg [33-1:0] _mystream_a30_source_count;
  reg [5-1:0] _mystream_a30_source_mode;
  reg [16-1:0] _mystream_a30_source_generator_id;
  reg [32-1:0] _mystream_a30_source_offset;
  reg [33-1:0] _mystream_a30_source_size;
  reg [32-1:0] _mystream_a30_source_stride;
  reg [32-1:0] _mystream_a30_source_offset_buf;
  reg [33-1:0] _mystream_a30_source_size_buf;
  reg [32-1:0] _mystream_a30_source_stride_buf;
  reg [8-1:0] _mystream_a30_source_sel;
  reg [32-1:0] _mystream_a30_source_ram_raddr;
  reg _mystream_a30_source_ram_renable;
  wire [32-1:0] _mystream_a30_source_ram_rdata;
  reg _mystream_a30_source_fifo_deq;
  wire [32-1:0] _mystream_a30_source_fifo_rdata;
  reg [32-1:0] _mystream_a30_source_empty_data;
  reg _mystream_a31_idle;
  reg [33-1:0] _mystream_a31_source_count;
  reg [5-1:0] _mystream_a31_source_mode;
  reg [16-1:0] _mystream_a31_source_generator_id;
  reg [32-1:0] _mystream_a31_source_offset;
  reg [33-1:0] _mystream_a31_source_size;
  reg [32-1:0] _mystream_a31_source_stride;
  reg [32-1:0] _mystream_a31_source_offset_buf;
  reg [33-1:0] _mystream_a31_source_size_buf;
  reg [32-1:0] _mystream_a31_source_stride_buf;
  reg [8-1:0] _mystream_a31_source_sel;
  reg [32-1:0] _mystream_a31_source_ram_raddr;
  reg _mystream_a31_source_ram_renable;
  wire [32-1:0] _mystream_a31_source_ram_rdata;
  reg _mystream_a31_source_fifo_deq;
  wire [32-1:0] _mystream_a31_source_fifo_rdata;
  reg [32-1:0] _mystream_a31_source_empty_data;
  reg _mystream_b0_idle;
  reg [33-1:0] _mystream_b0_source_count;
  reg [5-1:0] _mystream_b0_source_mode;
  reg [16-1:0] _mystream_b0_source_generator_id;
  reg [32-1:0] _mystream_b0_source_offset;
  reg [33-1:0] _mystream_b0_source_size;
  reg [32-1:0] _mystream_b0_source_stride;
  reg [32-1:0] _mystream_b0_source_offset_buf;
  reg [33-1:0] _mystream_b0_source_size_buf;
  reg [32-1:0] _mystream_b0_source_stride_buf;
  reg [8-1:0] _mystream_b0_source_sel;
  reg [32-1:0] _mystream_b0_source_ram_raddr;
  reg _mystream_b0_source_ram_renable;
  wire [32-1:0] _mystream_b0_source_ram_rdata;
  reg _mystream_b0_source_fifo_deq;
  wire [32-1:0] _mystream_b0_source_fifo_rdata;
  reg [32-1:0] _mystream_b0_source_empty_data;
  reg _mystream_b1_idle;
  reg [33-1:0] _mystream_b1_source_count;
  reg [5-1:0] _mystream_b1_source_mode;
  reg [16-1:0] _mystream_b1_source_generator_id;
  reg [32-1:0] _mystream_b1_source_offset;
  reg [33-1:0] _mystream_b1_source_size;
  reg [32-1:0] _mystream_b1_source_stride;
  reg [32-1:0] _mystream_b1_source_offset_buf;
  reg [33-1:0] _mystream_b1_source_size_buf;
  reg [32-1:0] _mystream_b1_source_stride_buf;
  reg [8-1:0] _mystream_b1_source_sel;
  reg [32-1:0] _mystream_b1_source_ram_raddr;
  reg _mystream_b1_source_ram_renable;
  wire [32-1:0] _mystream_b1_source_ram_rdata;
  reg _mystream_b1_source_fifo_deq;
  wire [32-1:0] _mystream_b1_source_fifo_rdata;
  reg [32-1:0] _mystream_b1_source_empty_data;
  reg _mystream_b2_idle;
  reg [33-1:0] _mystream_b2_source_count;
  reg [5-1:0] _mystream_b2_source_mode;
  reg [16-1:0] _mystream_b2_source_generator_id;
  reg [32-1:0] _mystream_b2_source_offset;
  reg [33-1:0] _mystream_b2_source_size;
  reg [32-1:0] _mystream_b2_source_stride;
  reg [32-1:0] _mystream_b2_source_offset_buf;
  reg [33-1:0] _mystream_b2_source_size_buf;
  reg [32-1:0] _mystream_b2_source_stride_buf;
  reg [8-1:0] _mystream_b2_source_sel;
  reg [32-1:0] _mystream_b2_source_ram_raddr;
  reg _mystream_b2_source_ram_renable;
  wire [32-1:0] _mystream_b2_source_ram_rdata;
  reg _mystream_b2_source_fifo_deq;
  wire [32-1:0] _mystream_b2_source_fifo_rdata;
  reg [32-1:0] _mystream_b2_source_empty_data;
  reg _mystream_b3_idle;
  reg [33-1:0] _mystream_b3_source_count;
  reg [5-1:0] _mystream_b3_source_mode;
  reg [16-1:0] _mystream_b3_source_generator_id;
  reg [32-1:0] _mystream_b3_source_offset;
  reg [33-1:0] _mystream_b3_source_size;
  reg [32-1:0] _mystream_b3_source_stride;
  reg [32-1:0] _mystream_b3_source_offset_buf;
  reg [33-1:0] _mystream_b3_source_size_buf;
  reg [32-1:0] _mystream_b3_source_stride_buf;
  reg [8-1:0] _mystream_b3_source_sel;
  reg [32-1:0] _mystream_b3_source_ram_raddr;
  reg _mystream_b3_source_ram_renable;
  wire [32-1:0] _mystream_b3_source_ram_rdata;
  reg _mystream_b3_source_fifo_deq;
  wire [32-1:0] _mystream_b3_source_fifo_rdata;
  reg [32-1:0] _mystream_b3_source_empty_data;
  reg _mystream_b4_idle;
  reg [33-1:0] _mystream_b4_source_count;
  reg [5-1:0] _mystream_b4_source_mode;
  reg [16-1:0] _mystream_b4_source_generator_id;
  reg [32-1:0] _mystream_b4_source_offset;
  reg [33-1:0] _mystream_b4_source_size;
  reg [32-1:0] _mystream_b4_source_stride;
  reg [32-1:0] _mystream_b4_source_offset_buf;
  reg [33-1:0] _mystream_b4_source_size_buf;
  reg [32-1:0] _mystream_b4_source_stride_buf;
  reg [8-1:0] _mystream_b4_source_sel;
  reg [32-1:0] _mystream_b4_source_ram_raddr;
  reg _mystream_b4_source_ram_renable;
  wire [32-1:0] _mystream_b4_source_ram_rdata;
  reg _mystream_b4_source_fifo_deq;
  wire [32-1:0] _mystream_b4_source_fifo_rdata;
  reg [32-1:0] _mystream_b4_source_empty_data;
  reg _mystream_b5_idle;
  reg [33-1:0] _mystream_b5_source_count;
  reg [5-1:0] _mystream_b5_source_mode;
  reg [16-1:0] _mystream_b5_source_generator_id;
  reg [32-1:0] _mystream_b5_source_offset;
  reg [33-1:0] _mystream_b5_source_size;
  reg [32-1:0] _mystream_b5_source_stride;
  reg [32-1:0] _mystream_b5_source_offset_buf;
  reg [33-1:0] _mystream_b5_source_size_buf;
  reg [32-1:0] _mystream_b5_source_stride_buf;
  reg [8-1:0] _mystream_b5_source_sel;
  reg [32-1:0] _mystream_b5_source_ram_raddr;
  reg _mystream_b5_source_ram_renable;
  wire [32-1:0] _mystream_b5_source_ram_rdata;
  reg _mystream_b5_source_fifo_deq;
  wire [32-1:0] _mystream_b5_source_fifo_rdata;
  reg [32-1:0] _mystream_b5_source_empty_data;
  reg _mystream_b6_idle;
  reg [33-1:0] _mystream_b6_source_count;
  reg [5-1:0] _mystream_b6_source_mode;
  reg [16-1:0] _mystream_b6_source_generator_id;
  reg [32-1:0] _mystream_b6_source_offset;
  reg [33-1:0] _mystream_b6_source_size;
  reg [32-1:0] _mystream_b6_source_stride;
  reg [32-1:0] _mystream_b6_source_offset_buf;
  reg [33-1:0] _mystream_b6_source_size_buf;
  reg [32-1:0] _mystream_b6_source_stride_buf;
  reg [8-1:0] _mystream_b6_source_sel;
  reg [32-1:0] _mystream_b6_source_ram_raddr;
  reg _mystream_b6_source_ram_renable;
  wire [32-1:0] _mystream_b6_source_ram_rdata;
  reg _mystream_b6_source_fifo_deq;
  wire [32-1:0] _mystream_b6_source_fifo_rdata;
  reg [32-1:0] _mystream_b6_source_empty_data;
  reg _mystream_b7_idle;
  reg [33-1:0] _mystream_b7_source_count;
  reg [5-1:0] _mystream_b7_source_mode;
  reg [16-1:0] _mystream_b7_source_generator_id;
  reg [32-1:0] _mystream_b7_source_offset;
  reg [33-1:0] _mystream_b7_source_size;
  reg [32-1:0] _mystream_b7_source_stride;
  reg [32-1:0] _mystream_b7_source_offset_buf;
  reg [33-1:0] _mystream_b7_source_size_buf;
  reg [32-1:0] _mystream_b7_source_stride_buf;
  reg [8-1:0] _mystream_b7_source_sel;
  reg [32-1:0] _mystream_b7_source_ram_raddr;
  reg _mystream_b7_source_ram_renable;
  wire [32-1:0] _mystream_b7_source_ram_rdata;
  reg _mystream_b7_source_fifo_deq;
  wire [32-1:0] _mystream_b7_source_fifo_rdata;
  reg [32-1:0] _mystream_b7_source_empty_data;
  reg _mystream_b8_idle;
  reg [33-1:0] _mystream_b8_source_count;
  reg [5-1:0] _mystream_b8_source_mode;
  reg [16-1:0] _mystream_b8_source_generator_id;
  reg [32-1:0] _mystream_b8_source_offset;
  reg [33-1:0] _mystream_b8_source_size;
  reg [32-1:0] _mystream_b8_source_stride;
  reg [32-1:0] _mystream_b8_source_offset_buf;
  reg [33-1:0] _mystream_b8_source_size_buf;
  reg [32-1:0] _mystream_b8_source_stride_buf;
  reg [8-1:0] _mystream_b8_source_sel;
  reg [32-1:0] _mystream_b8_source_ram_raddr;
  reg _mystream_b8_source_ram_renable;
  wire [32-1:0] _mystream_b8_source_ram_rdata;
  reg _mystream_b8_source_fifo_deq;
  wire [32-1:0] _mystream_b8_source_fifo_rdata;
  reg [32-1:0] _mystream_b8_source_empty_data;
  reg _mystream_b9_idle;
  reg [33-1:0] _mystream_b9_source_count;
  reg [5-1:0] _mystream_b9_source_mode;
  reg [16-1:0] _mystream_b9_source_generator_id;
  reg [32-1:0] _mystream_b9_source_offset;
  reg [33-1:0] _mystream_b9_source_size;
  reg [32-1:0] _mystream_b9_source_stride;
  reg [32-1:0] _mystream_b9_source_offset_buf;
  reg [33-1:0] _mystream_b9_source_size_buf;
  reg [32-1:0] _mystream_b9_source_stride_buf;
  reg [8-1:0] _mystream_b9_source_sel;
  reg [32-1:0] _mystream_b9_source_ram_raddr;
  reg _mystream_b9_source_ram_renable;
  wire [32-1:0] _mystream_b9_source_ram_rdata;
  reg _mystream_b9_source_fifo_deq;
  wire [32-1:0] _mystream_b9_source_fifo_rdata;
  reg [32-1:0] _mystream_b9_source_empty_data;
  reg _mystream_b10_idle;
  reg [33-1:0] _mystream_b10_source_count;
  reg [5-1:0] _mystream_b10_source_mode;
  reg [16-1:0] _mystream_b10_source_generator_id;
  reg [32-1:0] _mystream_b10_source_offset;
  reg [33-1:0] _mystream_b10_source_size;
  reg [32-1:0] _mystream_b10_source_stride;
  reg [32-1:0] _mystream_b10_source_offset_buf;
  reg [33-1:0] _mystream_b10_source_size_buf;
  reg [32-1:0] _mystream_b10_source_stride_buf;
  reg [8-1:0] _mystream_b10_source_sel;
  reg [32-1:0] _mystream_b10_source_ram_raddr;
  reg _mystream_b10_source_ram_renable;
  wire [32-1:0] _mystream_b10_source_ram_rdata;
  reg _mystream_b10_source_fifo_deq;
  wire [32-1:0] _mystream_b10_source_fifo_rdata;
  reg [32-1:0] _mystream_b10_source_empty_data;
  reg _mystream_b11_idle;
  reg [33-1:0] _mystream_b11_source_count;
  reg [5-1:0] _mystream_b11_source_mode;
  reg [16-1:0] _mystream_b11_source_generator_id;
  reg [32-1:0] _mystream_b11_source_offset;
  reg [33-1:0] _mystream_b11_source_size;
  reg [32-1:0] _mystream_b11_source_stride;
  reg [32-1:0] _mystream_b11_source_offset_buf;
  reg [33-1:0] _mystream_b11_source_size_buf;
  reg [32-1:0] _mystream_b11_source_stride_buf;
  reg [8-1:0] _mystream_b11_source_sel;
  reg [32-1:0] _mystream_b11_source_ram_raddr;
  reg _mystream_b11_source_ram_renable;
  wire [32-1:0] _mystream_b11_source_ram_rdata;
  reg _mystream_b11_source_fifo_deq;
  wire [32-1:0] _mystream_b11_source_fifo_rdata;
  reg [32-1:0] _mystream_b11_source_empty_data;
  reg _mystream_b12_idle;
  reg [33-1:0] _mystream_b12_source_count;
  reg [5-1:0] _mystream_b12_source_mode;
  reg [16-1:0] _mystream_b12_source_generator_id;
  reg [32-1:0] _mystream_b12_source_offset;
  reg [33-1:0] _mystream_b12_source_size;
  reg [32-1:0] _mystream_b12_source_stride;
  reg [32-1:0] _mystream_b12_source_offset_buf;
  reg [33-1:0] _mystream_b12_source_size_buf;
  reg [32-1:0] _mystream_b12_source_stride_buf;
  reg [8-1:0] _mystream_b12_source_sel;
  reg [32-1:0] _mystream_b12_source_ram_raddr;
  reg _mystream_b12_source_ram_renable;
  wire [32-1:0] _mystream_b12_source_ram_rdata;
  reg _mystream_b12_source_fifo_deq;
  wire [32-1:0] _mystream_b12_source_fifo_rdata;
  reg [32-1:0] _mystream_b12_source_empty_data;
  reg _mystream_b13_idle;
  reg [33-1:0] _mystream_b13_source_count;
  reg [5-1:0] _mystream_b13_source_mode;
  reg [16-1:0] _mystream_b13_source_generator_id;
  reg [32-1:0] _mystream_b13_source_offset;
  reg [33-1:0] _mystream_b13_source_size;
  reg [32-1:0] _mystream_b13_source_stride;
  reg [32-1:0] _mystream_b13_source_offset_buf;
  reg [33-1:0] _mystream_b13_source_size_buf;
  reg [32-1:0] _mystream_b13_source_stride_buf;
  reg [8-1:0] _mystream_b13_source_sel;
  reg [32-1:0] _mystream_b13_source_ram_raddr;
  reg _mystream_b13_source_ram_renable;
  wire [32-1:0] _mystream_b13_source_ram_rdata;
  reg _mystream_b13_source_fifo_deq;
  wire [32-1:0] _mystream_b13_source_fifo_rdata;
  reg [32-1:0] _mystream_b13_source_empty_data;
  reg _mystream_b14_idle;
  reg [33-1:0] _mystream_b14_source_count;
  reg [5-1:0] _mystream_b14_source_mode;
  reg [16-1:0] _mystream_b14_source_generator_id;
  reg [32-1:0] _mystream_b14_source_offset;
  reg [33-1:0] _mystream_b14_source_size;
  reg [32-1:0] _mystream_b14_source_stride;
  reg [32-1:0] _mystream_b14_source_offset_buf;
  reg [33-1:0] _mystream_b14_source_size_buf;
  reg [32-1:0] _mystream_b14_source_stride_buf;
  reg [8-1:0] _mystream_b14_source_sel;
  reg [32-1:0] _mystream_b14_source_ram_raddr;
  reg _mystream_b14_source_ram_renable;
  wire [32-1:0] _mystream_b14_source_ram_rdata;
  reg _mystream_b14_source_fifo_deq;
  wire [32-1:0] _mystream_b14_source_fifo_rdata;
  reg [32-1:0] _mystream_b14_source_empty_data;
  reg _mystream_b15_idle;
  reg [33-1:0] _mystream_b15_source_count;
  reg [5-1:0] _mystream_b15_source_mode;
  reg [16-1:0] _mystream_b15_source_generator_id;
  reg [32-1:0] _mystream_b15_source_offset;
  reg [33-1:0] _mystream_b15_source_size;
  reg [32-1:0] _mystream_b15_source_stride;
  reg [32-1:0] _mystream_b15_source_offset_buf;
  reg [33-1:0] _mystream_b15_source_size_buf;
  reg [32-1:0] _mystream_b15_source_stride_buf;
  reg [8-1:0] _mystream_b15_source_sel;
  reg [32-1:0] _mystream_b15_source_ram_raddr;
  reg _mystream_b15_source_ram_renable;
  wire [32-1:0] _mystream_b15_source_ram_rdata;
  reg _mystream_b15_source_fifo_deq;
  wire [32-1:0] _mystream_b15_source_fifo_rdata;
  reg [32-1:0] _mystream_b15_source_empty_data;
  reg _mystream_b16_idle;
  reg [33-1:0] _mystream_b16_source_count;
  reg [5-1:0] _mystream_b16_source_mode;
  reg [16-1:0] _mystream_b16_source_generator_id;
  reg [32-1:0] _mystream_b16_source_offset;
  reg [33-1:0] _mystream_b16_source_size;
  reg [32-1:0] _mystream_b16_source_stride;
  reg [32-1:0] _mystream_b16_source_offset_buf;
  reg [33-1:0] _mystream_b16_source_size_buf;
  reg [32-1:0] _mystream_b16_source_stride_buf;
  reg [8-1:0] _mystream_b16_source_sel;
  reg [32-1:0] _mystream_b16_source_ram_raddr;
  reg _mystream_b16_source_ram_renable;
  wire [32-1:0] _mystream_b16_source_ram_rdata;
  reg _mystream_b16_source_fifo_deq;
  wire [32-1:0] _mystream_b16_source_fifo_rdata;
  reg [32-1:0] _mystream_b16_source_empty_data;
  reg _mystream_b17_idle;
  reg [33-1:0] _mystream_b17_source_count;
  reg [5-1:0] _mystream_b17_source_mode;
  reg [16-1:0] _mystream_b17_source_generator_id;
  reg [32-1:0] _mystream_b17_source_offset;
  reg [33-1:0] _mystream_b17_source_size;
  reg [32-1:0] _mystream_b17_source_stride;
  reg [32-1:0] _mystream_b17_source_offset_buf;
  reg [33-1:0] _mystream_b17_source_size_buf;
  reg [32-1:0] _mystream_b17_source_stride_buf;
  reg [8-1:0] _mystream_b17_source_sel;
  reg [32-1:0] _mystream_b17_source_ram_raddr;
  reg _mystream_b17_source_ram_renable;
  wire [32-1:0] _mystream_b17_source_ram_rdata;
  reg _mystream_b17_source_fifo_deq;
  wire [32-1:0] _mystream_b17_source_fifo_rdata;
  reg [32-1:0] _mystream_b17_source_empty_data;
  reg _mystream_b18_idle;
  reg [33-1:0] _mystream_b18_source_count;
  reg [5-1:0] _mystream_b18_source_mode;
  reg [16-1:0] _mystream_b18_source_generator_id;
  reg [32-1:0] _mystream_b18_source_offset;
  reg [33-1:0] _mystream_b18_source_size;
  reg [32-1:0] _mystream_b18_source_stride;
  reg [32-1:0] _mystream_b18_source_offset_buf;
  reg [33-1:0] _mystream_b18_source_size_buf;
  reg [32-1:0] _mystream_b18_source_stride_buf;
  reg [8-1:0] _mystream_b18_source_sel;
  reg [32-1:0] _mystream_b18_source_ram_raddr;
  reg _mystream_b18_source_ram_renable;
  wire [32-1:0] _mystream_b18_source_ram_rdata;
  reg _mystream_b18_source_fifo_deq;
  wire [32-1:0] _mystream_b18_source_fifo_rdata;
  reg [32-1:0] _mystream_b18_source_empty_data;
  reg _mystream_b19_idle;
  reg [33-1:0] _mystream_b19_source_count;
  reg [5-1:0] _mystream_b19_source_mode;
  reg [16-1:0] _mystream_b19_source_generator_id;
  reg [32-1:0] _mystream_b19_source_offset;
  reg [33-1:0] _mystream_b19_source_size;
  reg [32-1:0] _mystream_b19_source_stride;
  reg [32-1:0] _mystream_b19_source_offset_buf;
  reg [33-1:0] _mystream_b19_source_size_buf;
  reg [32-1:0] _mystream_b19_source_stride_buf;
  reg [8-1:0] _mystream_b19_source_sel;
  reg [32-1:0] _mystream_b19_source_ram_raddr;
  reg _mystream_b19_source_ram_renable;
  wire [32-1:0] _mystream_b19_source_ram_rdata;
  reg _mystream_b19_source_fifo_deq;
  wire [32-1:0] _mystream_b19_source_fifo_rdata;
  reg [32-1:0] _mystream_b19_source_empty_data;
  reg _mystream_b20_idle;
  reg [33-1:0] _mystream_b20_source_count;
  reg [5-1:0] _mystream_b20_source_mode;
  reg [16-1:0] _mystream_b20_source_generator_id;
  reg [32-1:0] _mystream_b20_source_offset;
  reg [33-1:0] _mystream_b20_source_size;
  reg [32-1:0] _mystream_b20_source_stride;
  reg [32-1:0] _mystream_b20_source_offset_buf;
  reg [33-1:0] _mystream_b20_source_size_buf;
  reg [32-1:0] _mystream_b20_source_stride_buf;
  reg [8-1:0] _mystream_b20_source_sel;
  reg [32-1:0] _mystream_b20_source_ram_raddr;
  reg _mystream_b20_source_ram_renable;
  wire [32-1:0] _mystream_b20_source_ram_rdata;
  reg _mystream_b20_source_fifo_deq;
  wire [32-1:0] _mystream_b20_source_fifo_rdata;
  reg [32-1:0] _mystream_b20_source_empty_data;
  reg _mystream_b21_idle;
  reg [33-1:0] _mystream_b21_source_count;
  reg [5-1:0] _mystream_b21_source_mode;
  reg [16-1:0] _mystream_b21_source_generator_id;
  reg [32-1:0] _mystream_b21_source_offset;
  reg [33-1:0] _mystream_b21_source_size;
  reg [32-1:0] _mystream_b21_source_stride;
  reg [32-1:0] _mystream_b21_source_offset_buf;
  reg [33-1:0] _mystream_b21_source_size_buf;
  reg [32-1:0] _mystream_b21_source_stride_buf;
  reg [8-1:0] _mystream_b21_source_sel;
  reg [32-1:0] _mystream_b21_source_ram_raddr;
  reg _mystream_b21_source_ram_renable;
  wire [32-1:0] _mystream_b21_source_ram_rdata;
  reg _mystream_b21_source_fifo_deq;
  wire [32-1:0] _mystream_b21_source_fifo_rdata;
  reg [32-1:0] _mystream_b21_source_empty_data;
  reg _mystream_b22_idle;
  reg [33-1:0] _mystream_b22_source_count;
  reg [5-1:0] _mystream_b22_source_mode;
  reg [16-1:0] _mystream_b22_source_generator_id;
  reg [32-1:0] _mystream_b22_source_offset;
  reg [33-1:0] _mystream_b22_source_size;
  reg [32-1:0] _mystream_b22_source_stride;
  reg [32-1:0] _mystream_b22_source_offset_buf;
  reg [33-1:0] _mystream_b22_source_size_buf;
  reg [32-1:0] _mystream_b22_source_stride_buf;
  reg [8-1:0] _mystream_b22_source_sel;
  reg [32-1:0] _mystream_b22_source_ram_raddr;
  reg _mystream_b22_source_ram_renable;
  wire [32-1:0] _mystream_b22_source_ram_rdata;
  reg _mystream_b22_source_fifo_deq;
  wire [32-1:0] _mystream_b22_source_fifo_rdata;
  reg [32-1:0] _mystream_b22_source_empty_data;
  reg _mystream_b23_idle;
  reg [33-1:0] _mystream_b23_source_count;
  reg [5-1:0] _mystream_b23_source_mode;
  reg [16-1:0] _mystream_b23_source_generator_id;
  reg [32-1:0] _mystream_b23_source_offset;
  reg [33-1:0] _mystream_b23_source_size;
  reg [32-1:0] _mystream_b23_source_stride;
  reg [32-1:0] _mystream_b23_source_offset_buf;
  reg [33-1:0] _mystream_b23_source_size_buf;
  reg [32-1:0] _mystream_b23_source_stride_buf;
  reg [8-1:0] _mystream_b23_source_sel;
  reg [32-1:0] _mystream_b23_source_ram_raddr;
  reg _mystream_b23_source_ram_renable;
  wire [32-1:0] _mystream_b23_source_ram_rdata;
  reg _mystream_b23_source_fifo_deq;
  wire [32-1:0] _mystream_b23_source_fifo_rdata;
  reg [32-1:0] _mystream_b23_source_empty_data;
  reg _mystream_b24_idle;
  reg [33-1:0] _mystream_b24_source_count;
  reg [5-1:0] _mystream_b24_source_mode;
  reg [16-1:0] _mystream_b24_source_generator_id;
  reg [32-1:0] _mystream_b24_source_offset;
  reg [33-1:0] _mystream_b24_source_size;
  reg [32-1:0] _mystream_b24_source_stride;
  reg [32-1:0] _mystream_b24_source_offset_buf;
  reg [33-1:0] _mystream_b24_source_size_buf;
  reg [32-1:0] _mystream_b24_source_stride_buf;
  reg [8-1:0] _mystream_b24_source_sel;
  reg [32-1:0] _mystream_b24_source_ram_raddr;
  reg _mystream_b24_source_ram_renable;
  wire [32-1:0] _mystream_b24_source_ram_rdata;
  reg _mystream_b24_source_fifo_deq;
  wire [32-1:0] _mystream_b24_source_fifo_rdata;
  reg [32-1:0] _mystream_b24_source_empty_data;
  reg _mystream_b25_idle;
  reg [33-1:0] _mystream_b25_source_count;
  reg [5-1:0] _mystream_b25_source_mode;
  reg [16-1:0] _mystream_b25_source_generator_id;
  reg [32-1:0] _mystream_b25_source_offset;
  reg [33-1:0] _mystream_b25_source_size;
  reg [32-1:0] _mystream_b25_source_stride;
  reg [32-1:0] _mystream_b25_source_offset_buf;
  reg [33-1:0] _mystream_b25_source_size_buf;
  reg [32-1:0] _mystream_b25_source_stride_buf;
  reg [8-1:0] _mystream_b25_source_sel;
  reg [32-1:0] _mystream_b25_source_ram_raddr;
  reg _mystream_b25_source_ram_renable;
  wire [32-1:0] _mystream_b25_source_ram_rdata;
  reg _mystream_b25_source_fifo_deq;
  wire [32-1:0] _mystream_b25_source_fifo_rdata;
  reg [32-1:0] _mystream_b25_source_empty_data;
  reg _mystream_b26_idle;
  reg [33-1:0] _mystream_b26_source_count;
  reg [5-1:0] _mystream_b26_source_mode;
  reg [16-1:0] _mystream_b26_source_generator_id;
  reg [32-1:0] _mystream_b26_source_offset;
  reg [33-1:0] _mystream_b26_source_size;
  reg [32-1:0] _mystream_b26_source_stride;
  reg [32-1:0] _mystream_b26_source_offset_buf;
  reg [33-1:0] _mystream_b26_source_size_buf;
  reg [32-1:0] _mystream_b26_source_stride_buf;
  reg [8-1:0] _mystream_b26_source_sel;
  reg [32-1:0] _mystream_b26_source_ram_raddr;
  reg _mystream_b26_source_ram_renable;
  wire [32-1:0] _mystream_b26_source_ram_rdata;
  reg _mystream_b26_source_fifo_deq;
  wire [32-1:0] _mystream_b26_source_fifo_rdata;
  reg [32-1:0] _mystream_b26_source_empty_data;
  reg _mystream_b27_idle;
  reg [33-1:0] _mystream_b27_source_count;
  reg [5-1:0] _mystream_b27_source_mode;
  reg [16-1:0] _mystream_b27_source_generator_id;
  reg [32-1:0] _mystream_b27_source_offset;
  reg [33-1:0] _mystream_b27_source_size;
  reg [32-1:0] _mystream_b27_source_stride;
  reg [32-1:0] _mystream_b27_source_offset_buf;
  reg [33-1:0] _mystream_b27_source_size_buf;
  reg [32-1:0] _mystream_b27_source_stride_buf;
  reg [8-1:0] _mystream_b27_source_sel;
  reg [32-1:0] _mystream_b27_source_ram_raddr;
  reg _mystream_b27_source_ram_renable;
  wire [32-1:0] _mystream_b27_source_ram_rdata;
  reg _mystream_b27_source_fifo_deq;
  wire [32-1:0] _mystream_b27_source_fifo_rdata;
  reg [32-1:0] _mystream_b27_source_empty_data;
  reg _mystream_b28_idle;
  reg [33-1:0] _mystream_b28_source_count;
  reg [5-1:0] _mystream_b28_source_mode;
  reg [16-1:0] _mystream_b28_source_generator_id;
  reg [32-1:0] _mystream_b28_source_offset;
  reg [33-1:0] _mystream_b28_source_size;
  reg [32-1:0] _mystream_b28_source_stride;
  reg [32-1:0] _mystream_b28_source_offset_buf;
  reg [33-1:0] _mystream_b28_source_size_buf;
  reg [32-1:0] _mystream_b28_source_stride_buf;
  reg [8-1:0] _mystream_b28_source_sel;
  reg [32-1:0] _mystream_b28_source_ram_raddr;
  reg _mystream_b28_source_ram_renable;
  wire [32-1:0] _mystream_b28_source_ram_rdata;
  reg _mystream_b28_source_fifo_deq;
  wire [32-1:0] _mystream_b28_source_fifo_rdata;
  reg [32-1:0] _mystream_b28_source_empty_data;
  reg _mystream_b29_idle;
  reg [33-1:0] _mystream_b29_source_count;
  reg [5-1:0] _mystream_b29_source_mode;
  reg [16-1:0] _mystream_b29_source_generator_id;
  reg [32-1:0] _mystream_b29_source_offset;
  reg [33-1:0] _mystream_b29_source_size;
  reg [32-1:0] _mystream_b29_source_stride;
  reg [32-1:0] _mystream_b29_source_offset_buf;
  reg [33-1:0] _mystream_b29_source_size_buf;
  reg [32-1:0] _mystream_b29_source_stride_buf;
  reg [8-1:0] _mystream_b29_source_sel;
  reg [32-1:0] _mystream_b29_source_ram_raddr;
  reg _mystream_b29_source_ram_renable;
  wire [32-1:0] _mystream_b29_source_ram_rdata;
  reg _mystream_b29_source_fifo_deq;
  wire [32-1:0] _mystream_b29_source_fifo_rdata;
  reg [32-1:0] _mystream_b29_source_empty_data;
  reg _mystream_b30_idle;
  reg [33-1:0] _mystream_b30_source_count;
  reg [5-1:0] _mystream_b30_source_mode;
  reg [16-1:0] _mystream_b30_source_generator_id;
  reg [32-1:0] _mystream_b30_source_offset;
  reg [33-1:0] _mystream_b30_source_size;
  reg [32-1:0] _mystream_b30_source_stride;
  reg [32-1:0] _mystream_b30_source_offset_buf;
  reg [33-1:0] _mystream_b30_source_size_buf;
  reg [32-1:0] _mystream_b30_source_stride_buf;
  reg [8-1:0] _mystream_b30_source_sel;
  reg [32-1:0] _mystream_b30_source_ram_raddr;
  reg _mystream_b30_source_ram_renable;
  wire [32-1:0] _mystream_b30_source_ram_rdata;
  reg _mystream_b30_source_fifo_deq;
  wire [32-1:0] _mystream_b30_source_fifo_rdata;
  reg [32-1:0] _mystream_b30_source_empty_data;
  reg _mystream_b31_idle;
  reg [33-1:0] _mystream_b31_source_count;
  reg [5-1:0] _mystream_b31_source_mode;
  reg [16-1:0] _mystream_b31_source_generator_id;
  reg [32-1:0] _mystream_b31_source_offset;
  reg [33-1:0] _mystream_b31_source_size;
  reg [32-1:0] _mystream_b31_source_stride;
  reg [32-1:0] _mystream_b31_source_offset_buf;
  reg [33-1:0] _mystream_b31_source_size_buf;
  reg [32-1:0] _mystream_b31_source_stride_buf;
  reg [8-1:0] _mystream_b31_source_sel;
  reg [32-1:0] _mystream_b31_source_ram_raddr;
  reg _mystream_b31_source_ram_renable;
  wire [32-1:0] _mystream_b31_source_ram_rdata;
  reg _mystream_b31_source_fifo_deq;
  wire [32-1:0] _mystream_b31_source_fifo_rdata;
  reg [32-1:0] _mystream_b31_source_empty_data;
  reg _mystream_bias0_idle;
  reg [33-1:0] _mystream_bias0_source_count;
  reg [5-1:0] _mystream_bias0_source_mode;
  reg [16-1:0] _mystream_bias0_source_generator_id;
  reg [32-1:0] _mystream_bias0_source_offset;
  reg [33-1:0] _mystream_bias0_source_size;
  reg [32-1:0] _mystream_bias0_source_stride;
  reg [32-1:0] _mystream_bias0_source_offset_buf;
  reg [33-1:0] _mystream_bias0_source_size_buf;
  reg [32-1:0] _mystream_bias0_source_stride_buf;
  reg [8-1:0] _mystream_bias0_source_sel;
  reg [32-1:0] _mystream_bias0_source_ram_raddr;
  reg _mystream_bias0_source_ram_renable;
  wire [32-1:0] _mystream_bias0_source_ram_rdata;
  reg _mystream_bias0_source_fifo_deq;
  wire [32-1:0] _mystream_bias0_source_fifo_rdata;
  reg [32-1:0] _mystream_bias0_source_empty_data;
  reg _mystream_bias1_idle;
  reg [33-1:0] _mystream_bias1_source_count;
  reg [5-1:0] _mystream_bias1_source_mode;
  reg [16-1:0] _mystream_bias1_source_generator_id;
  reg [32-1:0] _mystream_bias1_source_offset;
  reg [33-1:0] _mystream_bias1_source_size;
  reg [32-1:0] _mystream_bias1_source_stride;
  reg [32-1:0] _mystream_bias1_source_offset_buf;
  reg [33-1:0] _mystream_bias1_source_size_buf;
  reg [32-1:0] _mystream_bias1_source_stride_buf;
  reg [8-1:0] _mystream_bias1_source_sel;
  reg [32-1:0] _mystream_bias1_source_ram_raddr;
  reg _mystream_bias1_source_ram_renable;
  wire [32-1:0] _mystream_bias1_source_ram_rdata;
  reg _mystream_bias1_source_fifo_deq;
  wire [32-1:0] _mystream_bias1_source_fifo_rdata;
  reg [32-1:0] _mystream_bias1_source_empty_data;
  reg _mystream_bias2_idle;
  reg [33-1:0] _mystream_bias2_source_count;
  reg [5-1:0] _mystream_bias2_source_mode;
  reg [16-1:0] _mystream_bias2_source_generator_id;
  reg [32-1:0] _mystream_bias2_source_offset;
  reg [33-1:0] _mystream_bias2_source_size;
  reg [32-1:0] _mystream_bias2_source_stride;
  reg [32-1:0] _mystream_bias2_source_offset_buf;
  reg [33-1:0] _mystream_bias2_source_size_buf;
  reg [32-1:0] _mystream_bias2_source_stride_buf;
  reg [8-1:0] _mystream_bias2_source_sel;
  reg [32-1:0] _mystream_bias2_source_ram_raddr;
  reg _mystream_bias2_source_ram_renable;
  wire [32-1:0] _mystream_bias2_source_ram_rdata;
  reg _mystream_bias2_source_fifo_deq;
  wire [32-1:0] _mystream_bias2_source_fifo_rdata;
  reg [32-1:0] _mystream_bias2_source_empty_data;
  reg _mystream_bias3_idle;
  reg [33-1:0] _mystream_bias3_source_count;
  reg [5-1:0] _mystream_bias3_source_mode;
  reg [16-1:0] _mystream_bias3_source_generator_id;
  reg [32-1:0] _mystream_bias3_source_offset;
  reg [33-1:0] _mystream_bias3_source_size;
  reg [32-1:0] _mystream_bias3_source_stride;
  reg [32-1:0] _mystream_bias3_source_offset_buf;
  reg [33-1:0] _mystream_bias3_source_size_buf;
  reg [32-1:0] _mystream_bias3_source_stride_buf;
  reg [8-1:0] _mystream_bias3_source_sel;
  reg [32-1:0] _mystream_bias3_source_ram_raddr;
  reg _mystream_bias3_source_ram_renable;
  wire [32-1:0] _mystream_bias3_source_ram_rdata;
  reg _mystream_bias3_source_fifo_deq;
  wire [32-1:0] _mystream_bias3_source_fifo_rdata;
  reg [32-1:0] _mystream_bias3_source_empty_data;
  reg _mystream_bias4_idle;
  reg [33-1:0] _mystream_bias4_source_count;
  reg [5-1:0] _mystream_bias4_source_mode;
  reg [16-1:0] _mystream_bias4_source_generator_id;
  reg [32-1:0] _mystream_bias4_source_offset;
  reg [33-1:0] _mystream_bias4_source_size;
  reg [32-1:0] _mystream_bias4_source_stride;
  reg [32-1:0] _mystream_bias4_source_offset_buf;
  reg [33-1:0] _mystream_bias4_source_size_buf;
  reg [32-1:0] _mystream_bias4_source_stride_buf;
  reg [8-1:0] _mystream_bias4_source_sel;
  reg [32-1:0] _mystream_bias4_source_ram_raddr;
  reg _mystream_bias4_source_ram_renable;
  wire [32-1:0] _mystream_bias4_source_ram_rdata;
  reg _mystream_bias4_source_fifo_deq;
  wire [32-1:0] _mystream_bias4_source_fifo_rdata;
  reg [32-1:0] _mystream_bias4_source_empty_data;
  reg _mystream_bias5_idle;
  reg [33-1:0] _mystream_bias5_source_count;
  reg [5-1:0] _mystream_bias5_source_mode;
  reg [16-1:0] _mystream_bias5_source_generator_id;
  reg [32-1:0] _mystream_bias5_source_offset;
  reg [33-1:0] _mystream_bias5_source_size;
  reg [32-1:0] _mystream_bias5_source_stride;
  reg [32-1:0] _mystream_bias5_source_offset_buf;
  reg [33-1:0] _mystream_bias5_source_size_buf;
  reg [32-1:0] _mystream_bias5_source_stride_buf;
  reg [8-1:0] _mystream_bias5_source_sel;
  reg [32-1:0] _mystream_bias5_source_ram_raddr;
  reg _mystream_bias5_source_ram_renable;
  wire [32-1:0] _mystream_bias5_source_ram_rdata;
  reg _mystream_bias5_source_fifo_deq;
  wire [32-1:0] _mystream_bias5_source_fifo_rdata;
  reg [32-1:0] _mystream_bias5_source_empty_data;
  reg _mystream_bias6_idle;
  reg [33-1:0] _mystream_bias6_source_count;
  reg [5-1:0] _mystream_bias6_source_mode;
  reg [16-1:0] _mystream_bias6_source_generator_id;
  reg [32-1:0] _mystream_bias6_source_offset;
  reg [33-1:0] _mystream_bias6_source_size;
  reg [32-1:0] _mystream_bias6_source_stride;
  reg [32-1:0] _mystream_bias6_source_offset_buf;
  reg [33-1:0] _mystream_bias6_source_size_buf;
  reg [32-1:0] _mystream_bias6_source_stride_buf;
  reg [8-1:0] _mystream_bias6_source_sel;
  reg [32-1:0] _mystream_bias6_source_ram_raddr;
  reg _mystream_bias6_source_ram_renable;
  wire [32-1:0] _mystream_bias6_source_ram_rdata;
  reg _mystream_bias6_source_fifo_deq;
  wire [32-1:0] _mystream_bias6_source_fifo_rdata;
  reg [32-1:0] _mystream_bias6_source_empty_data;
  reg _mystream_bias7_idle;
  reg [33-1:0] _mystream_bias7_source_count;
  reg [5-1:0] _mystream_bias7_source_mode;
  reg [16-1:0] _mystream_bias7_source_generator_id;
  reg [32-1:0] _mystream_bias7_source_offset;
  reg [33-1:0] _mystream_bias7_source_size;
  reg [32-1:0] _mystream_bias7_source_stride;
  reg [32-1:0] _mystream_bias7_source_offset_buf;
  reg [33-1:0] _mystream_bias7_source_size_buf;
  reg [32-1:0] _mystream_bias7_source_stride_buf;
  reg [8-1:0] _mystream_bias7_source_sel;
  reg [32-1:0] _mystream_bias7_source_ram_raddr;
  reg _mystream_bias7_source_ram_renable;
  wire [32-1:0] _mystream_bias7_source_ram_rdata;
  reg _mystream_bias7_source_fifo_deq;
  wire [32-1:0] _mystream_bias7_source_fifo_rdata;
  reg [32-1:0] _mystream_bias7_source_empty_data;
  reg _mystream_bias8_idle;
  reg [33-1:0] _mystream_bias8_source_count;
  reg [5-1:0] _mystream_bias8_source_mode;
  reg [16-1:0] _mystream_bias8_source_generator_id;
  reg [32-1:0] _mystream_bias8_source_offset;
  reg [33-1:0] _mystream_bias8_source_size;
  reg [32-1:0] _mystream_bias8_source_stride;
  reg [32-1:0] _mystream_bias8_source_offset_buf;
  reg [33-1:0] _mystream_bias8_source_size_buf;
  reg [32-1:0] _mystream_bias8_source_stride_buf;
  reg [8-1:0] _mystream_bias8_source_sel;
  reg [32-1:0] _mystream_bias8_source_ram_raddr;
  reg _mystream_bias8_source_ram_renable;
  wire [32-1:0] _mystream_bias8_source_ram_rdata;
  reg _mystream_bias8_source_fifo_deq;
  wire [32-1:0] _mystream_bias8_source_fifo_rdata;
  reg [32-1:0] _mystream_bias8_source_empty_data;
  reg _mystream_bias9_idle;
  reg [33-1:0] _mystream_bias9_source_count;
  reg [5-1:0] _mystream_bias9_source_mode;
  reg [16-1:0] _mystream_bias9_source_generator_id;
  reg [32-1:0] _mystream_bias9_source_offset;
  reg [33-1:0] _mystream_bias9_source_size;
  reg [32-1:0] _mystream_bias9_source_stride;
  reg [32-1:0] _mystream_bias9_source_offset_buf;
  reg [33-1:0] _mystream_bias9_source_size_buf;
  reg [32-1:0] _mystream_bias9_source_stride_buf;
  reg [8-1:0] _mystream_bias9_source_sel;
  reg [32-1:0] _mystream_bias9_source_ram_raddr;
  reg _mystream_bias9_source_ram_renable;
  wire [32-1:0] _mystream_bias9_source_ram_rdata;
  reg _mystream_bias9_source_fifo_deq;
  wire [32-1:0] _mystream_bias9_source_fifo_rdata;
  reg [32-1:0] _mystream_bias9_source_empty_data;
  reg _mystream_bias10_idle;
  reg [33-1:0] _mystream_bias10_source_count;
  reg [5-1:0] _mystream_bias10_source_mode;
  reg [16-1:0] _mystream_bias10_source_generator_id;
  reg [32-1:0] _mystream_bias10_source_offset;
  reg [33-1:0] _mystream_bias10_source_size;
  reg [32-1:0] _mystream_bias10_source_stride;
  reg [32-1:0] _mystream_bias10_source_offset_buf;
  reg [33-1:0] _mystream_bias10_source_size_buf;
  reg [32-1:0] _mystream_bias10_source_stride_buf;
  reg [8-1:0] _mystream_bias10_source_sel;
  reg [32-1:0] _mystream_bias10_source_ram_raddr;
  reg _mystream_bias10_source_ram_renable;
  wire [32-1:0] _mystream_bias10_source_ram_rdata;
  reg _mystream_bias10_source_fifo_deq;
  wire [32-1:0] _mystream_bias10_source_fifo_rdata;
  reg [32-1:0] _mystream_bias10_source_empty_data;
  reg _mystream_bias11_idle;
  reg [33-1:0] _mystream_bias11_source_count;
  reg [5-1:0] _mystream_bias11_source_mode;
  reg [16-1:0] _mystream_bias11_source_generator_id;
  reg [32-1:0] _mystream_bias11_source_offset;
  reg [33-1:0] _mystream_bias11_source_size;
  reg [32-1:0] _mystream_bias11_source_stride;
  reg [32-1:0] _mystream_bias11_source_offset_buf;
  reg [33-1:0] _mystream_bias11_source_size_buf;
  reg [32-1:0] _mystream_bias11_source_stride_buf;
  reg [8-1:0] _mystream_bias11_source_sel;
  reg [32-1:0] _mystream_bias11_source_ram_raddr;
  reg _mystream_bias11_source_ram_renable;
  wire [32-1:0] _mystream_bias11_source_ram_rdata;
  reg _mystream_bias11_source_fifo_deq;
  wire [32-1:0] _mystream_bias11_source_fifo_rdata;
  reg [32-1:0] _mystream_bias11_source_empty_data;
  reg _mystream_bias12_idle;
  reg [33-1:0] _mystream_bias12_source_count;
  reg [5-1:0] _mystream_bias12_source_mode;
  reg [16-1:0] _mystream_bias12_source_generator_id;
  reg [32-1:0] _mystream_bias12_source_offset;
  reg [33-1:0] _mystream_bias12_source_size;
  reg [32-1:0] _mystream_bias12_source_stride;
  reg [32-1:0] _mystream_bias12_source_offset_buf;
  reg [33-1:0] _mystream_bias12_source_size_buf;
  reg [32-1:0] _mystream_bias12_source_stride_buf;
  reg [8-1:0] _mystream_bias12_source_sel;
  reg [32-1:0] _mystream_bias12_source_ram_raddr;
  reg _mystream_bias12_source_ram_renable;
  wire [32-1:0] _mystream_bias12_source_ram_rdata;
  reg _mystream_bias12_source_fifo_deq;
  wire [32-1:0] _mystream_bias12_source_fifo_rdata;
  reg [32-1:0] _mystream_bias12_source_empty_data;
  reg _mystream_bias13_idle;
  reg [33-1:0] _mystream_bias13_source_count;
  reg [5-1:0] _mystream_bias13_source_mode;
  reg [16-1:0] _mystream_bias13_source_generator_id;
  reg [32-1:0] _mystream_bias13_source_offset;
  reg [33-1:0] _mystream_bias13_source_size;
  reg [32-1:0] _mystream_bias13_source_stride;
  reg [32-1:0] _mystream_bias13_source_offset_buf;
  reg [33-1:0] _mystream_bias13_source_size_buf;
  reg [32-1:0] _mystream_bias13_source_stride_buf;
  reg [8-1:0] _mystream_bias13_source_sel;
  reg [32-1:0] _mystream_bias13_source_ram_raddr;
  reg _mystream_bias13_source_ram_renable;
  wire [32-1:0] _mystream_bias13_source_ram_rdata;
  reg _mystream_bias13_source_fifo_deq;
  wire [32-1:0] _mystream_bias13_source_fifo_rdata;
  reg [32-1:0] _mystream_bias13_source_empty_data;
  reg _mystream_bias14_idle;
  reg [33-1:0] _mystream_bias14_source_count;
  reg [5-1:0] _mystream_bias14_source_mode;
  reg [16-1:0] _mystream_bias14_source_generator_id;
  reg [32-1:0] _mystream_bias14_source_offset;
  reg [33-1:0] _mystream_bias14_source_size;
  reg [32-1:0] _mystream_bias14_source_stride;
  reg [32-1:0] _mystream_bias14_source_offset_buf;
  reg [33-1:0] _mystream_bias14_source_size_buf;
  reg [32-1:0] _mystream_bias14_source_stride_buf;
  reg [8-1:0] _mystream_bias14_source_sel;
  reg [32-1:0] _mystream_bias14_source_ram_raddr;
  reg _mystream_bias14_source_ram_renable;
  wire [32-1:0] _mystream_bias14_source_ram_rdata;
  reg _mystream_bias14_source_fifo_deq;
  wire [32-1:0] _mystream_bias14_source_fifo_rdata;
  reg [32-1:0] _mystream_bias14_source_empty_data;
  reg _mystream_bias15_idle;
  reg [33-1:0] _mystream_bias15_source_count;
  reg [5-1:0] _mystream_bias15_source_mode;
  reg [16-1:0] _mystream_bias15_source_generator_id;
  reg [32-1:0] _mystream_bias15_source_offset;
  reg [33-1:0] _mystream_bias15_source_size;
  reg [32-1:0] _mystream_bias15_source_stride;
  reg [32-1:0] _mystream_bias15_source_offset_buf;
  reg [33-1:0] _mystream_bias15_source_size_buf;
  reg [32-1:0] _mystream_bias15_source_stride_buf;
  reg [8-1:0] _mystream_bias15_source_sel;
  reg [32-1:0] _mystream_bias15_source_ram_raddr;
  reg _mystream_bias15_source_ram_renable;
  wire [32-1:0] _mystream_bias15_source_ram_rdata;
  reg _mystream_bias15_source_fifo_deq;
  wire [32-1:0] _mystream_bias15_source_fifo_rdata;
  reg [32-1:0] _mystream_bias15_source_empty_data;
  reg _mystream_bias16_idle;
  reg [33-1:0] _mystream_bias16_source_count;
  reg [5-1:0] _mystream_bias16_source_mode;
  reg [16-1:0] _mystream_bias16_source_generator_id;
  reg [32-1:0] _mystream_bias16_source_offset;
  reg [33-1:0] _mystream_bias16_source_size;
  reg [32-1:0] _mystream_bias16_source_stride;
  reg [32-1:0] _mystream_bias16_source_offset_buf;
  reg [33-1:0] _mystream_bias16_source_size_buf;
  reg [32-1:0] _mystream_bias16_source_stride_buf;
  reg [8-1:0] _mystream_bias16_source_sel;
  reg [32-1:0] _mystream_bias16_source_ram_raddr;
  reg _mystream_bias16_source_ram_renable;
  wire [32-1:0] _mystream_bias16_source_ram_rdata;
  reg _mystream_bias16_source_fifo_deq;
  wire [32-1:0] _mystream_bias16_source_fifo_rdata;
  reg [32-1:0] _mystream_bias16_source_empty_data;
  reg _mystream_bias17_idle;
  reg [33-1:0] _mystream_bias17_source_count;
  reg [5-1:0] _mystream_bias17_source_mode;
  reg [16-1:0] _mystream_bias17_source_generator_id;
  reg [32-1:0] _mystream_bias17_source_offset;
  reg [33-1:0] _mystream_bias17_source_size;
  reg [32-1:0] _mystream_bias17_source_stride;
  reg [32-1:0] _mystream_bias17_source_offset_buf;
  reg [33-1:0] _mystream_bias17_source_size_buf;
  reg [32-1:0] _mystream_bias17_source_stride_buf;
  reg [8-1:0] _mystream_bias17_source_sel;
  reg [32-1:0] _mystream_bias17_source_ram_raddr;
  reg _mystream_bias17_source_ram_renable;
  wire [32-1:0] _mystream_bias17_source_ram_rdata;
  reg _mystream_bias17_source_fifo_deq;
  wire [32-1:0] _mystream_bias17_source_fifo_rdata;
  reg [32-1:0] _mystream_bias17_source_empty_data;
  reg _mystream_bias18_idle;
  reg [33-1:0] _mystream_bias18_source_count;
  reg [5-1:0] _mystream_bias18_source_mode;
  reg [16-1:0] _mystream_bias18_source_generator_id;
  reg [32-1:0] _mystream_bias18_source_offset;
  reg [33-1:0] _mystream_bias18_source_size;
  reg [32-1:0] _mystream_bias18_source_stride;
  reg [32-1:0] _mystream_bias18_source_offset_buf;
  reg [33-1:0] _mystream_bias18_source_size_buf;
  reg [32-1:0] _mystream_bias18_source_stride_buf;
  reg [8-1:0] _mystream_bias18_source_sel;
  reg [32-1:0] _mystream_bias18_source_ram_raddr;
  reg _mystream_bias18_source_ram_renable;
  wire [32-1:0] _mystream_bias18_source_ram_rdata;
  reg _mystream_bias18_source_fifo_deq;
  wire [32-1:0] _mystream_bias18_source_fifo_rdata;
  reg [32-1:0] _mystream_bias18_source_empty_data;
  reg _mystream_bias19_idle;
  reg [33-1:0] _mystream_bias19_source_count;
  reg [5-1:0] _mystream_bias19_source_mode;
  reg [16-1:0] _mystream_bias19_source_generator_id;
  reg [32-1:0] _mystream_bias19_source_offset;
  reg [33-1:0] _mystream_bias19_source_size;
  reg [32-1:0] _mystream_bias19_source_stride;
  reg [32-1:0] _mystream_bias19_source_offset_buf;
  reg [33-1:0] _mystream_bias19_source_size_buf;
  reg [32-1:0] _mystream_bias19_source_stride_buf;
  reg [8-1:0] _mystream_bias19_source_sel;
  reg [32-1:0] _mystream_bias19_source_ram_raddr;
  reg _mystream_bias19_source_ram_renable;
  wire [32-1:0] _mystream_bias19_source_ram_rdata;
  reg _mystream_bias19_source_fifo_deq;
  wire [32-1:0] _mystream_bias19_source_fifo_rdata;
  reg [32-1:0] _mystream_bias19_source_empty_data;
  reg _mystream_bias20_idle;
  reg [33-1:0] _mystream_bias20_source_count;
  reg [5-1:0] _mystream_bias20_source_mode;
  reg [16-1:0] _mystream_bias20_source_generator_id;
  reg [32-1:0] _mystream_bias20_source_offset;
  reg [33-1:0] _mystream_bias20_source_size;
  reg [32-1:0] _mystream_bias20_source_stride;
  reg [32-1:0] _mystream_bias20_source_offset_buf;
  reg [33-1:0] _mystream_bias20_source_size_buf;
  reg [32-1:0] _mystream_bias20_source_stride_buf;
  reg [8-1:0] _mystream_bias20_source_sel;
  reg [32-1:0] _mystream_bias20_source_ram_raddr;
  reg _mystream_bias20_source_ram_renable;
  wire [32-1:0] _mystream_bias20_source_ram_rdata;
  reg _mystream_bias20_source_fifo_deq;
  wire [32-1:0] _mystream_bias20_source_fifo_rdata;
  reg [32-1:0] _mystream_bias20_source_empty_data;
  reg _mystream_bias21_idle;
  reg [33-1:0] _mystream_bias21_source_count;
  reg [5-1:0] _mystream_bias21_source_mode;
  reg [16-1:0] _mystream_bias21_source_generator_id;
  reg [32-1:0] _mystream_bias21_source_offset;
  reg [33-1:0] _mystream_bias21_source_size;
  reg [32-1:0] _mystream_bias21_source_stride;
  reg [32-1:0] _mystream_bias21_source_offset_buf;
  reg [33-1:0] _mystream_bias21_source_size_buf;
  reg [32-1:0] _mystream_bias21_source_stride_buf;
  reg [8-1:0] _mystream_bias21_source_sel;
  reg [32-1:0] _mystream_bias21_source_ram_raddr;
  reg _mystream_bias21_source_ram_renable;
  wire [32-1:0] _mystream_bias21_source_ram_rdata;
  reg _mystream_bias21_source_fifo_deq;
  wire [32-1:0] _mystream_bias21_source_fifo_rdata;
  reg [32-1:0] _mystream_bias21_source_empty_data;
  reg _mystream_bias22_idle;
  reg [33-1:0] _mystream_bias22_source_count;
  reg [5-1:0] _mystream_bias22_source_mode;
  reg [16-1:0] _mystream_bias22_source_generator_id;
  reg [32-1:0] _mystream_bias22_source_offset;
  reg [33-1:0] _mystream_bias22_source_size;
  reg [32-1:0] _mystream_bias22_source_stride;
  reg [32-1:0] _mystream_bias22_source_offset_buf;
  reg [33-1:0] _mystream_bias22_source_size_buf;
  reg [32-1:0] _mystream_bias22_source_stride_buf;
  reg [8-1:0] _mystream_bias22_source_sel;
  reg [32-1:0] _mystream_bias22_source_ram_raddr;
  reg _mystream_bias22_source_ram_renable;
  wire [32-1:0] _mystream_bias22_source_ram_rdata;
  reg _mystream_bias22_source_fifo_deq;
  wire [32-1:0] _mystream_bias22_source_fifo_rdata;
  reg [32-1:0] _mystream_bias22_source_empty_data;
  reg _mystream_bias23_idle;
  reg [33-1:0] _mystream_bias23_source_count;
  reg [5-1:0] _mystream_bias23_source_mode;
  reg [16-1:0] _mystream_bias23_source_generator_id;
  reg [32-1:0] _mystream_bias23_source_offset;
  reg [33-1:0] _mystream_bias23_source_size;
  reg [32-1:0] _mystream_bias23_source_stride;
  reg [32-1:0] _mystream_bias23_source_offset_buf;
  reg [33-1:0] _mystream_bias23_source_size_buf;
  reg [32-1:0] _mystream_bias23_source_stride_buf;
  reg [8-1:0] _mystream_bias23_source_sel;
  reg [32-1:0] _mystream_bias23_source_ram_raddr;
  reg _mystream_bias23_source_ram_renable;
  wire [32-1:0] _mystream_bias23_source_ram_rdata;
  reg _mystream_bias23_source_fifo_deq;
  wire [32-1:0] _mystream_bias23_source_fifo_rdata;
  reg [32-1:0] _mystream_bias23_source_empty_data;
  reg _mystream_bias24_idle;
  reg [33-1:0] _mystream_bias24_source_count;
  reg [5-1:0] _mystream_bias24_source_mode;
  reg [16-1:0] _mystream_bias24_source_generator_id;
  reg [32-1:0] _mystream_bias24_source_offset;
  reg [33-1:0] _mystream_bias24_source_size;
  reg [32-1:0] _mystream_bias24_source_stride;
  reg [32-1:0] _mystream_bias24_source_offset_buf;
  reg [33-1:0] _mystream_bias24_source_size_buf;
  reg [32-1:0] _mystream_bias24_source_stride_buf;
  reg [8-1:0] _mystream_bias24_source_sel;
  reg [32-1:0] _mystream_bias24_source_ram_raddr;
  reg _mystream_bias24_source_ram_renable;
  wire [32-1:0] _mystream_bias24_source_ram_rdata;
  reg _mystream_bias24_source_fifo_deq;
  wire [32-1:0] _mystream_bias24_source_fifo_rdata;
  reg [32-1:0] _mystream_bias24_source_empty_data;
  reg _mystream_bias25_idle;
  reg [33-1:0] _mystream_bias25_source_count;
  reg [5-1:0] _mystream_bias25_source_mode;
  reg [16-1:0] _mystream_bias25_source_generator_id;
  reg [32-1:0] _mystream_bias25_source_offset;
  reg [33-1:0] _mystream_bias25_source_size;
  reg [32-1:0] _mystream_bias25_source_stride;
  reg [32-1:0] _mystream_bias25_source_offset_buf;
  reg [33-1:0] _mystream_bias25_source_size_buf;
  reg [32-1:0] _mystream_bias25_source_stride_buf;
  reg [8-1:0] _mystream_bias25_source_sel;
  reg [32-1:0] _mystream_bias25_source_ram_raddr;
  reg _mystream_bias25_source_ram_renable;
  wire [32-1:0] _mystream_bias25_source_ram_rdata;
  reg _mystream_bias25_source_fifo_deq;
  wire [32-1:0] _mystream_bias25_source_fifo_rdata;
  reg [32-1:0] _mystream_bias25_source_empty_data;
  reg _mystream_bias26_idle;
  reg [33-1:0] _mystream_bias26_source_count;
  reg [5-1:0] _mystream_bias26_source_mode;
  reg [16-1:0] _mystream_bias26_source_generator_id;
  reg [32-1:0] _mystream_bias26_source_offset;
  reg [33-1:0] _mystream_bias26_source_size;
  reg [32-1:0] _mystream_bias26_source_stride;
  reg [32-1:0] _mystream_bias26_source_offset_buf;
  reg [33-1:0] _mystream_bias26_source_size_buf;
  reg [32-1:0] _mystream_bias26_source_stride_buf;
  reg [8-1:0] _mystream_bias26_source_sel;
  reg [32-1:0] _mystream_bias26_source_ram_raddr;
  reg _mystream_bias26_source_ram_renable;
  wire [32-1:0] _mystream_bias26_source_ram_rdata;
  reg _mystream_bias26_source_fifo_deq;
  wire [32-1:0] _mystream_bias26_source_fifo_rdata;
  reg [32-1:0] _mystream_bias26_source_empty_data;
  reg _mystream_bias27_idle;
  reg [33-1:0] _mystream_bias27_source_count;
  reg [5-1:0] _mystream_bias27_source_mode;
  reg [16-1:0] _mystream_bias27_source_generator_id;
  reg [32-1:0] _mystream_bias27_source_offset;
  reg [33-1:0] _mystream_bias27_source_size;
  reg [32-1:0] _mystream_bias27_source_stride;
  reg [32-1:0] _mystream_bias27_source_offset_buf;
  reg [33-1:0] _mystream_bias27_source_size_buf;
  reg [32-1:0] _mystream_bias27_source_stride_buf;
  reg [8-1:0] _mystream_bias27_source_sel;
  reg [32-1:0] _mystream_bias27_source_ram_raddr;
  reg _mystream_bias27_source_ram_renable;
  wire [32-1:0] _mystream_bias27_source_ram_rdata;
  reg _mystream_bias27_source_fifo_deq;
  wire [32-1:0] _mystream_bias27_source_fifo_rdata;
  reg [32-1:0] _mystream_bias27_source_empty_data;
  reg _mystream_bias28_idle;
  reg [33-1:0] _mystream_bias28_source_count;
  reg [5-1:0] _mystream_bias28_source_mode;
  reg [16-1:0] _mystream_bias28_source_generator_id;
  reg [32-1:0] _mystream_bias28_source_offset;
  reg [33-1:0] _mystream_bias28_source_size;
  reg [32-1:0] _mystream_bias28_source_stride;
  reg [32-1:0] _mystream_bias28_source_offset_buf;
  reg [33-1:0] _mystream_bias28_source_size_buf;
  reg [32-1:0] _mystream_bias28_source_stride_buf;
  reg [8-1:0] _mystream_bias28_source_sel;
  reg [32-1:0] _mystream_bias28_source_ram_raddr;
  reg _mystream_bias28_source_ram_renable;
  wire [32-1:0] _mystream_bias28_source_ram_rdata;
  reg _mystream_bias28_source_fifo_deq;
  wire [32-1:0] _mystream_bias28_source_fifo_rdata;
  reg [32-1:0] _mystream_bias28_source_empty_data;
  reg _mystream_bias29_idle;
  reg [33-1:0] _mystream_bias29_source_count;
  reg [5-1:0] _mystream_bias29_source_mode;
  reg [16-1:0] _mystream_bias29_source_generator_id;
  reg [32-1:0] _mystream_bias29_source_offset;
  reg [33-1:0] _mystream_bias29_source_size;
  reg [32-1:0] _mystream_bias29_source_stride;
  reg [32-1:0] _mystream_bias29_source_offset_buf;
  reg [33-1:0] _mystream_bias29_source_size_buf;
  reg [32-1:0] _mystream_bias29_source_stride_buf;
  reg [8-1:0] _mystream_bias29_source_sel;
  reg [32-1:0] _mystream_bias29_source_ram_raddr;
  reg _mystream_bias29_source_ram_renable;
  wire [32-1:0] _mystream_bias29_source_ram_rdata;
  reg _mystream_bias29_source_fifo_deq;
  wire [32-1:0] _mystream_bias29_source_fifo_rdata;
  reg [32-1:0] _mystream_bias29_source_empty_data;
  reg _mystream_bias30_idle;
  reg [33-1:0] _mystream_bias30_source_count;
  reg [5-1:0] _mystream_bias30_source_mode;
  reg [16-1:0] _mystream_bias30_source_generator_id;
  reg [32-1:0] _mystream_bias30_source_offset;
  reg [33-1:0] _mystream_bias30_source_size;
  reg [32-1:0] _mystream_bias30_source_stride;
  reg [32-1:0] _mystream_bias30_source_offset_buf;
  reg [33-1:0] _mystream_bias30_source_size_buf;
  reg [32-1:0] _mystream_bias30_source_stride_buf;
  reg [8-1:0] _mystream_bias30_source_sel;
  reg [32-1:0] _mystream_bias30_source_ram_raddr;
  reg _mystream_bias30_source_ram_renable;
  wire [32-1:0] _mystream_bias30_source_ram_rdata;
  reg _mystream_bias30_source_fifo_deq;
  wire [32-1:0] _mystream_bias30_source_fifo_rdata;
  reg [32-1:0] _mystream_bias30_source_empty_data;
  reg _mystream_bias31_idle;
  reg [33-1:0] _mystream_bias31_source_count;
  reg [5-1:0] _mystream_bias31_source_mode;
  reg [16-1:0] _mystream_bias31_source_generator_id;
  reg [32-1:0] _mystream_bias31_source_offset;
  reg [33-1:0] _mystream_bias31_source_size;
  reg [32-1:0] _mystream_bias31_source_stride;
  reg [32-1:0] _mystream_bias31_source_offset_buf;
  reg [33-1:0] _mystream_bias31_source_size_buf;
  reg [32-1:0] _mystream_bias31_source_stride_buf;
  reg [8-1:0] _mystream_bias31_source_sel;
  reg [32-1:0] _mystream_bias31_source_ram_raddr;
  reg _mystream_bias31_source_ram_renable;
  wire [32-1:0] _mystream_bias31_source_ram_rdata;
  reg _mystream_bias31_source_fifo_deq;
  wire [32-1:0] _mystream_bias31_source_fifo_rdata;
  reg [32-1:0] _mystream_bias31_source_empty_data;
  reg [33-1:0] _mystream_sum_vec0_sink_count;
  reg [5-1:0] _mystream_sum_vec0_sink_mode;
  reg [16-1:0] _mystream_sum_vec0_sink_generator_id;
  reg [32-1:0] _mystream_sum_vec0_sink_offset;
  reg [33-1:0] _mystream_sum_vec0_sink_size;
  reg [32-1:0] _mystream_sum_vec0_sink_stride;
  reg [32-1:0] _mystream_sum_vec0_sink_offset_buf;
  reg [33-1:0] _mystream_sum_vec0_sink_size_buf;
  reg [32-1:0] _mystream_sum_vec0_sink_stride_buf;
  reg [8-1:0] _mystream_sum_vec0_sink_sel;
  reg [32-1:0] _mystream_sum_vec0_sink_waddr;
  reg _mystream_sum_vec0_sink_wenable;
  reg [32-1:0] _mystream_sum_vec0_sink_wdata;
  reg _mystream_sum_vec0_sink_fifo_enq;
  reg [32-1:0] _mystream_sum_vec0_sink_fifo_wdata;
  reg [32-1:0] _mystream_sum_vec0_sink_immediate;
  reg [33-1:0] _mystream_sum_vec1_sink_count;
  reg [5-1:0] _mystream_sum_vec1_sink_mode;
  reg [16-1:0] _mystream_sum_vec1_sink_generator_id;
  reg [32-1:0] _mystream_sum_vec1_sink_offset;
  reg [33-1:0] _mystream_sum_vec1_sink_size;
  reg [32-1:0] _mystream_sum_vec1_sink_stride;
  reg [32-1:0] _mystream_sum_vec1_sink_offset_buf;
  reg [33-1:0] _mystream_sum_vec1_sink_size_buf;
  reg [32-1:0] _mystream_sum_vec1_sink_stride_buf;
  reg [8-1:0] _mystream_sum_vec1_sink_sel;
  reg [32-1:0] _mystream_sum_vec1_sink_waddr;
  reg _mystream_sum_vec1_sink_wenable;
  reg [32-1:0] _mystream_sum_vec1_sink_wdata;
  reg _mystream_sum_vec1_sink_fifo_enq;
  reg [32-1:0] _mystream_sum_vec1_sink_fifo_wdata;
  reg [32-1:0] _mystream_sum_vec1_sink_immediate;
  reg [33-1:0] _mystream_sum_vec2_sink_count;
  reg [5-1:0] _mystream_sum_vec2_sink_mode;
  reg [16-1:0] _mystream_sum_vec2_sink_generator_id;
  reg [32-1:0] _mystream_sum_vec2_sink_offset;
  reg [33-1:0] _mystream_sum_vec2_sink_size;
  reg [32-1:0] _mystream_sum_vec2_sink_stride;
  reg [32-1:0] _mystream_sum_vec2_sink_offset_buf;
  reg [33-1:0] _mystream_sum_vec2_sink_size_buf;
  reg [32-1:0] _mystream_sum_vec2_sink_stride_buf;
  reg [8-1:0] _mystream_sum_vec2_sink_sel;
  reg [32-1:0] _mystream_sum_vec2_sink_waddr;
  reg _mystream_sum_vec2_sink_wenable;
  reg [32-1:0] _mystream_sum_vec2_sink_wdata;
  reg _mystream_sum_vec2_sink_fifo_enq;
  reg [32-1:0] _mystream_sum_vec2_sink_fifo_wdata;
  reg [32-1:0] _mystream_sum_vec2_sink_immediate;
  reg [33-1:0] _mystream_sum_vec3_sink_count;
  reg [5-1:0] _mystream_sum_vec3_sink_mode;
  reg [16-1:0] _mystream_sum_vec3_sink_generator_id;
  reg [32-1:0] _mystream_sum_vec3_sink_offset;
  reg [33-1:0] _mystream_sum_vec3_sink_size;
  reg [32-1:0] _mystream_sum_vec3_sink_stride;
  reg [32-1:0] _mystream_sum_vec3_sink_offset_buf;
  reg [33-1:0] _mystream_sum_vec3_sink_size_buf;
  reg [32-1:0] _mystream_sum_vec3_sink_stride_buf;
  reg [8-1:0] _mystream_sum_vec3_sink_sel;
  reg [32-1:0] _mystream_sum_vec3_sink_waddr;
  reg _mystream_sum_vec3_sink_wenable;
  reg [32-1:0] _mystream_sum_vec3_sink_wdata;
  reg _mystream_sum_vec3_sink_fifo_enq;
  reg [32-1:0] _mystream_sum_vec3_sink_fifo_wdata;
  reg [32-1:0] _mystream_sum_vec3_sink_immediate;
  reg [33-1:0] _mystream_sum_vec4_sink_count;
  reg [5-1:0] _mystream_sum_vec4_sink_mode;
  reg [16-1:0] _mystream_sum_vec4_sink_generator_id;
  reg [32-1:0] _mystream_sum_vec4_sink_offset;
  reg [33-1:0] _mystream_sum_vec4_sink_size;
  reg [32-1:0] _mystream_sum_vec4_sink_stride;
  reg [32-1:0] _mystream_sum_vec4_sink_offset_buf;
  reg [33-1:0] _mystream_sum_vec4_sink_size_buf;
  reg [32-1:0] _mystream_sum_vec4_sink_stride_buf;
  reg [8-1:0] _mystream_sum_vec4_sink_sel;
  reg [32-1:0] _mystream_sum_vec4_sink_waddr;
  reg _mystream_sum_vec4_sink_wenable;
  reg [32-1:0] _mystream_sum_vec4_sink_wdata;
  reg _mystream_sum_vec4_sink_fifo_enq;
  reg [32-1:0] _mystream_sum_vec4_sink_fifo_wdata;
  reg [32-1:0] _mystream_sum_vec4_sink_immediate;
  reg [33-1:0] _mystream_sum_vec5_sink_count;
  reg [5-1:0] _mystream_sum_vec5_sink_mode;
  reg [16-1:0] _mystream_sum_vec5_sink_generator_id;
  reg [32-1:0] _mystream_sum_vec5_sink_offset;
  reg [33-1:0] _mystream_sum_vec5_sink_size;
  reg [32-1:0] _mystream_sum_vec5_sink_stride;
  reg [32-1:0] _mystream_sum_vec5_sink_offset_buf;
  reg [33-1:0] _mystream_sum_vec5_sink_size_buf;
  reg [32-1:0] _mystream_sum_vec5_sink_stride_buf;
  reg [8-1:0] _mystream_sum_vec5_sink_sel;
  reg [32-1:0] _mystream_sum_vec5_sink_waddr;
  reg _mystream_sum_vec5_sink_wenable;
  reg [32-1:0] _mystream_sum_vec5_sink_wdata;
  reg _mystream_sum_vec5_sink_fifo_enq;
  reg [32-1:0] _mystream_sum_vec5_sink_fifo_wdata;
  reg [32-1:0] _mystream_sum_vec5_sink_immediate;
  reg [33-1:0] _mystream_sum_vec6_sink_count;
  reg [5-1:0] _mystream_sum_vec6_sink_mode;
  reg [16-1:0] _mystream_sum_vec6_sink_generator_id;
  reg [32-1:0] _mystream_sum_vec6_sink_offset;
  reg [33-1:0] _mystream_sum_vec6_sink_size;
  reg [32-1:0] _mystream_sum_vec6_sink_stride;
  reg [32-1:0] _mystream_sum_vec6_sink_offset_buf;
  reg [33-1:0] _mystream_sum_vec6_sink_size_buf;
  reg [32-1:0] _mystream_sum_vec6_sink_stride_buf;
  reg [8-1:0] _mystream_sum_vec6_sink_sel;
  reg [32-1:0] _mystream_sum_vec6_sink_waddr;
  reg _mystream_sum_vec6_sink_wenable;
  reg [32-1:0] _mystream_sum_vec6_sink_wdata;
  reg _mystream_sum_vec6_sink_fifo_enq;
  reg [32-1:0] _mystream_sum_vec6_sink_fifo_wdata;
  reg [32-1:0] _mystream_sum_vec6_sink_immediate;
  reg [33-1:0] _mystream_sum_vec7_sink_count;
  reg [5-1:0] _mystream_sum_vec7_sink_mode;
  reg [16-1:0] _mystream_sum_vec7_sink_generator_id;
  reg [32-1:0] _mystream_sum_vec7_sink_offset;
  reg [33-1:0] _mystream_sum_vec7_sink_size;
  reg [32-1:0] _mystream_sum_vec7_sink_stride;
  reg [32-1:0] _mystream_sum_vec7_sink_offset_buf;
  reg [33-1:0] _mystream_sum_vec7_sink_size_buf;
  reg [32-1:0] _mystream_sum_vec7_sink_stride_buf;
  reg [8-1:0] _mystream_sum_vec7_sink_sel;
  reg [32-1:0] _mystream_sum_vec7_sink_waddr;
  reg _mystream_sum_vec7_sink_wenable;
  reg [32-1:0] _mystream_sum_vec7_sink_wdata;
  reg _mystream_sum_vec7_sink_fifo_enq;
  reg [32-1:0] _mystream_sum_vec7_sink_fifo_wdata;
  reg [32-1:0] _mystream_sum_vec7_sink_immediate;
  reg [33-1:0] _mystream_sum_vec8_sink_count;
  reg [5-1:0] _mystream_sum_vec8_sink_mode;
  reg [16-1:0] _mystream_sum_vec8_sink_generator_id;
  reg [32-1:0] _mystream_sum_vec8_sink_offset;
  reg [33-1:0] _mystream_sum_vec8_sink_size;
  reg [32-1:0] _mystream_sum_vec8_sink_stride;
  reg [32-1:0] _mystream_sum_vec8_sink_offset_buf;
  reg [33-1:0] _mystream_sum_vec8_sink_size_buf;
  reg [32-1:0] _mystream_sum_vec8_sink_stride_buf;
  reg [8-1:0] _mystream_sum_vec8_sink_sel;
  reg [32-1:0] _mystream_sum_vec8_sink_waddr;
  reg _mystream_sum_vec8_sink_wenable;
  reg [32-1:0] _mystream_sum_vec8_sink_wdata;
  reg _mystream_sum_vec8_sink_fifo_enq;
  reg [32-1:0] _mystream_sum_vec8_sink_fifo_wdata;
  reg [32-1:0] _mystream_sum_vec8_sink_immediate;
  reg [33-1:0] _mystream_sum_vec9_sink_count;
  reg [5-1:0] _mystream_sum_vec9_sink_mode;
  reg [16-1:0] _mystream_sum_vec9_sink_generator_id;
  reg [32-1:0] _mystream_sum_vec9_sink_offset;
  reg [33-1:0] _mystream_sum_vec9_sink_size;
  reg [32-1:0] _mystream_sum_vec9_sink_stride;
  reg [32-1:0] _mystream_sum_vec9_sink_offset_buf;
  reg [33-1:0] _mystream_sum_vec9_sink_size_buf;
  reg [32-1:0] _mystream_sum_vec9_sink_stride_buf;
  reg [8-1:0] _mystream_sum_vec9_sink_sel;
  reg [32-1:0] _mystream_sum_vec9_sink_waddr;
  reg _mystream_sum_vec9_sink_wenable;
  reg [32-1:0] _mystream_sum_vec9_sink_wdata;
  reg _mystream_sum_vec9_sink_fifo_enq;
  reg [32-1:0] _mystream_sum_vec9_sink_fifo_wdata;
  reg [32-1:0] _mystream_sum_vec9_sink_immediate;
  reg [33-1:0] _mystream_sum_vec10_sink_count;
  reg [5-1:0] _mystream_sum_vec10_sink_mode;
  reg [16-1:0] _mystream_sum_vec10_sink_generator_id;
  reg [32-1:0] _mystream_sum_vec10_sink_offset;
  reg [33-1:0] _mystream_sum_vec10_sink_size;
  reg [32-1:0] _mystream_sum_vec10_sink_stride;
  reg [32-1:0] _mystream_sum_vec10_sink_offset_buf;
  reg [33-1:0] _mystream_sum_vec10_sink_size_buf;
  reg [32-1:0] _mystream_sum_vec10_sink_stride_buf;
  reg [8-1:0] _mystream_sum_vec10_sink_sel;
  reg [32-1:0] _mystream_sum_vec10_sink_waddr;
  reg _mystream_sum_vec10_sink_wenable;
  reg [32-1:0] _mystream_sum_vec10_sink_wdata;
  reg _mystream_sum_vec10_sink_fifo_enq;
  reg [32-1:0] _mystream_sum_vec10_sink_fifo_wdata;
  reg [32-1:0] _mystream_sum_vec10_sink_immediate;
  reg [33-1:0] _mystream_sum_vec11_sink_count;
  reg [5-1:0] _mystream_sum_vec11_sink_mode;
  reg [16-1:0] _mystream_sum_vec11_sink_generator_id;
  reg [32-1:0] _mystream_sum_vec11_sink_offset;
  reg [33-1:0] _mystream_sum_vec11_sink_size;
  reg [32-1:0] _mystream_sum_vec11_sink_stride;
  reg [32-1:0] _mystream_sum_vec11_sink_offset_buf;
  reg [33-1:0] _mystream_sum_vec11_sink_size_buf;
  reg [32-1:0] _mystream_sum_vec11_sink_stride_buf;
  reg [8-1:0] _mystream_sum_vec11_sink_sel;
  reg [32-1:0] _mystream_sum_vec11_sink_waddr;
  reg _mystream_sum_vec11_sink_wenable;
  reg [32-1:0] _mystream_sum_vec11_sink_wdata;
  reg _mystream_sum_vec11_sink_fifo_enq;
  reg [32-1:0] _mystream_sum_vec11_sink_fifo_wdata;
  reg [32-1:0] _mystream_sum_vec11_sink_immediate;
  reg [33-1:0] _mystream_sum_vec12_sink_count;
  reg [5-1:0] _mystream_sum_vec12_sink_mode;
  reg [16-1:0] _mystream_sum_vec12_sink_generator_id;
  reg [32-1:0] _mystream_sum_vec12_sink_offset;
  reg [33-1:0] _mystream_sum_vec12_sink_size;
  reg [32-1:0] _mystream_sum_vec12_sink_stride;
  reg [32-1:0] _mystream_sum_vec12_sink_offset_buf;
  reg [33-1:0] _mystream_sum_vec12_sink_size_buf;
  reg [32-1:0] _mystream_sum_vec12_sink_stride_buf;
  reg [8-1:0] _mystream_sum_vec12_sink_sel;
  reg [32-1:0] _mystream_sum_vec12_sink_waddr;
  reg _mystream_sum_vec12_sink_wenable;
  reg [32-1:0] _mystream_sum_vec12_sink_wdata;
  reg _mystream_sum_vec12_sink_fifo_enq;
  reg [32-1:0] _mystream_sum_vec12_sink_fifo_wdata;
  reg [32-1:0] _mystream_sum_vec12_sink_immediate;
  reg [33-1:0] _mystream_sum_vec13_sink_count;
  reg [5-1:0] _mystream_sum_vec13_sink_mode;
  reg [16-1:0] _mystream_sum_vec13_sink_generator_id;
  reg [32-1:0] _mystream_sum_vec13_sink_offset;
  reg [33-1:0] _mystream_sum_vec13_sink_size;
  reg [32-1:0] _mystream_sum_vec13_sink_stride;
  reg [32-1:0] _mystream_sum_vec13_sink_offset_buf;
  reg [33-1:0] _mystream_sum_vec13_sink_size_buf;
  reg [32-1:0] _mystream_sum_vec13_sink_stride_buf;
  reg [8-1:0] _mystream_sum_vec13_sink_sel;
  reg [32-1:0] _mystream_sum_vec13_sink_waddr;
  reg _mystream_sum_vec13_sink_wenable;
  reg [32-1:0] _mystream_sum_vec13_sink_wdata;
  reg _mystream_sum_vec13_sink_fifo_enq;
  reg [32-1:0] _mystream_sum_vec13_sink_fifo_wdata;
  reg [32-1:0] _mystream_sum_vec13_sink_immediate;
  reg [33-1:0] _mystream_sum_vec14_sink_count;
  reg [5-1:0] _mystream_sum_vec14_sink_mode;
  reg [16-1:0] _mystream_sum_vec14_sink_generator_id;
  reg [32-1:0] _mystream_sum_vec14_sink_offset;
  reg [33-1:0] _mystream_sum_vec14_sink_size;
  reg [32-1:0] _mystream_sum_vec14_sink_stride;
  reg [32-1:0] _mystream_sum_vec14_sink_offset_buf;
  reg [33-1:0] _mystream_sum_vec14_sink_size_buf;
  reg [32-1:0] _mystream_sum_vec14_sink_stride_buf;
  reg [8-1:0] _mystream_sum_vec14_sink_sel;
  reg [32-1:0] _mystream_sum_vec14_sink_waddr;
  reg _mystream_sum_vec14_sink_wenable;
  reg [32-1:0] _mystream_sum_vec14_sink_wdata;
  reg _mystream_sum_vec14_sink_fifo_enq;
  reg [32-1:0] _mystream_sum_vec14_sink_fifo_wdata;
  reg [32-1:0] _mystream_sum_vec14_sink_immediate;
  reg [33-1:0] _mystream_sum_vec15_sink_count;
  reg [5-1:0] _mystream_sum_vec15_sink_mode;
  reg [16-1:0] _mystream_sum_vec15_sink_generator_id;
  reg [32-1:0] _mystream_sum_vec15_sink_offset;
  reg [33-1:0] _mystream_sum_vec15_sink_size;
  reg [32-1:0] _mystream_sum_vec15_sink_stride;
  reg [32-1:0] _mystream_sum_vec15_sink_offset_buf;
  reg [33-1:0] _mystream_sum_vec15_sink_size_buf;
  reg [32-1:0] _mystream_sum_vec15_sink_stride_buf;
  reg [8-1:0] _mystream_sum_vec15_sink_sel;
  reg [32-1:0] _mystream_sum_vec15_sink_waddr;
  reg _mystream_sum_vec15_sink_wenable;
  reg [32-1:0] _mystream_sum_vec15_sink_wdata;
  reg _mystream_sum_vec15_sink_fifo_enq;
  reg [32-1:0] _mystream_sum_vec15_sink_fifo_wdata;
  reg [32-1:0] _mystream_sum_vec15_sink_immediate;
  reg [33-1:0] _mystream_sum_vec16_sink_count;
  reg [5-1:0] _mystream_sum_vec16_sink_mode;
  reg [16-1:0] _mystream_sum_vec16_sink_generator_id;
  reg [32-1:0] _mystream_sum_vec16_sink_offset;
  reg [33-1:0] _mystream_sum_vec16_sink_size;
  reg [32-1:0] _mystream_sum_vec16_sink_stride;
  reg [32-1:0] _mystream_sum_vec16_sink_offset_buf;
  reg [33-1:0] _mystream_sum_vec16_sink_size_buf;
  reg [32-1:0] _mystream_sum_vec16_sink_stride_buf;
  reg [8-1:0] _mystream_sum_vec16_sink_sel;
  reg [32-1:0] _mystream_sum_vec16_sink_waddr;
  reg _mystream_sum_vec16_sink_wenable;
  reg [32-1:0] _mystream_sum_vec16_sink_wdata;
  reg _mystream_sum_vec16_sink_fifo_enq;
  reg [32-1:0] _mystream_sum_vec16_sink_fifo_wdata;
  reg [32-1:0] _mystream_sum_vec16_sink_immediate;
  reg [33-1:0] _mystream_sum_vec17_sink_count;
  reg [5-1:0] _mystream_sum_vec17_sink_mode;
  reg [16-1:0] _mystream_sum_vec17_sink_generator_id;
  reg [32-1:0] _mystream_sum_vec17_sink_offset;
  reg [33-1:0] _mystream_sum_vec17_sink_size;
  reg [32-1:0] _mystream_sum_vec17_sink_stride;
  reg [32-1:0] _mystream_sum_vec17_sink_offset_buf;
  reg [33-1:0] _mystream_sum_vec17_sink_size_buf;
  reg [32-1:0] _mystream_sum_vec17_sink_stride_buf;
  reg [8-1:0] _mystream_sum_vec17_sink_sel;
  reg [32-1:0] _mystream_sum_vec17_sink_waddr;
  reg _mystream_sum_vec17_sink_wenable;
  reg [32-1:0] _mystream_sum_vec17_sink_wdata;
  reg _mystream_sum_vec17_sink_fifo_enq;
  reg [32-1:0] _mystream_sum_vec17_sink_fifo_wdata;
  reg [32-1:0] _mystream_sum_vec17_sink_immediate;
  reg [33-1:0] _mystream_sum_vec18_sink_count;
  reg [5-1:0] _mystream_sum_vec18_sink_mode;
  reg [16-1:0] _mystream_sum_vec18_sink_generator_id;
  reg [32-1:0] _mystream_sum_vec18_sink_offset;
  reg [33-1:0] _mystream_sum_vec18_sink_size;
  reg [32-1:0] _mystream_sum_vec18_sink_stride;
  reg [32-1:0] _mystream_sum_vec18_sink_offset_buf;
  reg [33-1:0] _mystream_sum_vec18_sink_size_buf;
  reg [32-1:0] _mystream_sum_vec18_sink_stride_buf;
  reg [8-1:0] _mystream_sum_vec18_sink_sel;
  reg [32-1:0] _mystream_sum_vec18_sink_waddr;
  reg _mystream_sum_vec18_sink_wenable;
  reg [32-1:0] _mystream_sum_vec18_sink_wdata;
  reg _mystream_sum_vec18_sink_fifo_enq;
  reg [32-1:0] _mystream_sum_vec18_sink_fifo_wdata;
  reg [32-1:0] _mystream_sum_vec18_sink_immediate;
  reg [33-1:0] _mystream_sum_vec19_sink_count;
  reg [5-1:0] _mystream_sum_vec19_sink_mode;
  reg [16-1:0] _mystream_sum_vec19_sink_generator_id;
  reg [32-1:0] _mystream_sum_vec19_sink_offset;
  reg [33-1:0] _mystream_sum_vec19_sink_size;
  reg [32-1:0] _mystream_sum_vec19_sink_stride;
  reg [32-1:0] _mystream_sum_vec19_sink_offset_buf;
  reg [33-1:0] _mystream_sum_vec19_sink_size_buf;
  reg [32-1:0] _mystream_sum_vec19_sink_stride_buf;
  reg [8-1:0] _mystream_sum_vec19_sink_sel;
  reg [32-1:0] _mystream_sum_vec19_sink_waddr;
  reg _mystream_sum_vec19_sink_wenable;
  reg [32-1:0] _mystream_sum_vec19_sink_wdata;
  reg _mystream_sum_vec19_sink_fifo_enq;
  reg [32-1:0] _mystream_sum_vec19_sink_fifo_wdata;
  reg [32-1:0] _mystream_sum_vec19_sink_immediate;
  reg [33-1:0] _mystream_sum_vec20_sink_count;
  reg [5-1:0] _mystream_sum_vec20_sink_mode;
  reg [16-1:0] _mystream_sum_vec20_sink_generator_id;
  reg [32-1:0] _mystream_sum_vec20_sink_offset;
  reg [33-1:0] _mystream_sum_vec20_sink_size;
  reg [32-1:0] _mystream_sum_vec20_sink_stride;
  reg [32-1:0] _mystream_sum_vec20_sink_offset_buf;
  reg [33-1:0] _mystream_sum_vec20_sink_size_buf;
  reg [32-1:0] _mystream_sum_vec20_sink_stride_buf;
  reg [8-1:0] _mystream_sum_vec20_sink_sel;
  reg [32-1:0] _mystream_sum_vec20_sink_waddr;
  reg _mystream_sum_vec20_sink_wenable;
  reg [32-1:0] _mystream_sum_vec20_sink_wdata;
  reg _mystream_sum_vec20_sink_fifo_enq;
  reg [32-1:0] _mystream_sum_vec20_sink_fifo_wdata;
  reg [32-1:0] _mystream_sum_vec20_sink_immediate;
  reg [33-1:0] _mystream_sum_vec21_sink_count;
  reg [5-1:0] _mystream_sum_vec21_sink_mode;
  reg [16-1:0] _mystream_sum_vec21_sink_generator_id;
  reg [32-1:0] _mystream_sum_vec21_sink_offset;
  reg [33-1:0] _mystream_sum_vec21_sink_size;
  reg [32-1:0] _mystream_sum_vec21_sink_stride;
  reg [32-1:0] _mystream_sum_vec21_sink_offset_buf;
  reg [33-1:0] _mystream_sum_vec21_sink_size_buf;
  reg [32-1:0] _mystream_sum_vec21_sink_stride_buf;
  reg [8-1:0] _mystream_sum_vec21_sink_sel;
  reg [32-1:0] _mystream_sum_vec21_sink_waddr;
  reg _mystream_sum_vec21_sink_wenable;
  reg [32-1:0] _mystream_sum_vec21_sink_wdata;
  reg _mystream_sum_vec21_sink_fifo_enq;
  reg [32-1:0] _mystream_sum_vec21_sink_fifo_wdata;
  reg [32-1:0] _mystream_sum_vec21_sink_immediate;
  reg [33-1:0] _mystream_sum_vec22_sink_count;
  reg [5-1:0] _mystream_sum_vec22_sink_mode;
  reg [16-1:0] _mystream_sum_vec22_sink_generator_id;
  reg [32-1:0] _mystream_sum_vec22_sink_offset;
  reg [33-1:0] _mystream_sum_vec22_sink_size;
  reg [32-1:0] _mystream_sum_vec22_sink_stride;
  reg [32-1:0] _mystream_sum_vec22_sink_offset_buf;
  reg [33-1:0] _mystream_sum_vec22_sink_size_buf;
  reg [32-1:0] _mystream_sum_vec22_sink_stride_buf;
  reg [8-1:0] _mystream_sum_vec22_sink_sel;
  reg [32-1:0] _mystream_sum_vec22_sink_waddr;
  reg _mystream_sum_vec22_sink_wenable;
  reg [32-1:0] _mystream_sum_vec22_sink_wdata;
  reg _mystream_sum_vec22_sink_fifo_enq;
  reg [32-1:0] _mystream_sum_vec22_sink_fifo_wdata;
  reg [32-1:0] _mystream_sum_vec22_sink_immediate;
  reg [33-1:0] _mystream_sum_vec23_sink_count;
  reg [5-1:0] _mystream_sum_vec23_sink_mode;
  reg [16-1:0] _mystream_sum_vec23_sink_generator_id;
  reg [32-1:0] _mystream_sum_vec23_sink_offset;
  reg [33-1:0] _mystream_sum_vec23_sink_size;
  reg [32-1:0] _mystream_sum_vec23_sink_stride;
  reg [32-1:0] _mystream_sum_vec23_sink_offset_buf;
  reg [33-1:0] _mystream_sum_vec23_sink_size_buf;
  reg [32-1:0] _mystream_sum_vec23_sink_stride_buf;
  reg [8-1:0] _mystream_sum_vec23_sink_sel;
  reg [32-1:0] _mystream_sum_vec23_sink_waddr;
  reg _mystream_sum_vec23_sink_wenable;
  reg [32-1:0] _mystream_sum_vec23_sink_wdata;
  reg _mystream_sum_vec23_sink_fifo_enq;
  reg [32-1:0] _mystream_sum_vec23_sink_fifo_wdata;
  reg [32-1:0] _mystream_sum_vec23_sink_immediate;
  reg [33-1:0] _mystream_sum_vec24_sink_count;
  reg [5-1:0] _mystream_sum_vec24_sink_mode;
  reg [16-1:0] _mystream_sum_vec24_sink_generator_id;
  reg [32-1:0] _mystream_sum_vec24_sink_offset;
  reg [33-1:0] _mystream_sum_vec24_sink_size;
  reg [32-1:0] _mystream_sum_vec24_sink_stride;
  reg [32-1:0] _mystream_sum_vec24_sink_offset_buf;
  reg [33-1:0] _mystream_sum_vec24_sink_size_buf;
  reg [32-1:0] _mystream_sum_vec24_sink_stride_buf;
  reg [8-1:0] _mystream_sum_vec24_sink_sel;
  reg [32-1:0] _mystream_sum_vec24_sink_waddr;
  reg _mystream_sum_vec24_sink_wenable;
  reg [32-1:0] _mystream_sum_vec24_sink_wdata;
  reg _mystream_sum_vec24_sink_fifo_enq;
  reg [32-1:0] _mystream_sum_vec24_sink_fifo_wdata;
  reg [32-1:0] _mystream_sum_vec24_sink_immediate;
  reg [33-1:0] _mystream_sum_vec25_sink_count;
  reg [5-1:0] _mystream_sum_vec25_sink_mode;
  reg [16-1:0] _mystream_sum_vec25_sink_generator_id;
  reg [32-1:0] _mystream_sum_vec25_sink_offset;
  reg [33-1:0] _mystream_sum_vec25_sink_size;
  reg [32-1:0] _mystream_sum_vec25_sink_stride;
  reg [32-1:0] _mystream_sum_vec25_sink_offset_buf;
  reg [33-1:0] _mystream_sum_vec25_sink_size_buf;
  reg [32-1:0] _mystream_sum_vec25_sink_stride_buf;
  reg [8-1:0] _mystream_sum_vec25_sink_sel;
  reg [32-1:0] _mystream_sum_vec25_sink_waddr;
  reg _mystream_sum_vec25_sink_wenable;
  reg [32-1:0] _mystream_sum_vec25_sink_wdata;
  reg _mystream_sum_vec25_sink_fifo_enq;
  reg [32-1:0] _mystream_sum_vec25_sink_fifo_wdata;
  reg [32-1:0] _mystream_sum_vec25_sink_immediate;
  reg [33-1:0] _mystream_sum_vec26_sink_count;
  reg [5-1:0] _mystream_sum_vec26_sink_mode;
  reg [16-1:0] _mystream_sum_vec26_sink_generator_id;
  reg [32-1:0] _mystream_sum_vec26_sink_offset;
  reg [33-1:0] _mystream_sum_vec26_sink_size;
  reg [32-1:0] _mystream_sum_vec26_sink_stride;
  reg [32-1:0] _mystream_sum_vec26_sink_offset_buf;
  reg [33-1:0] _mystream_sum_vec26_sink_size_buf;
  reg [32-1:0] _mystream_sum_vec26_sink_stride_buf;
  reg [8-1:0] _mystream_sum_vec26_sink_sel;
  reg [32-1:0] _mystream_sum_vec26_sink_waddr;
  reg _mystream_sum_vec26_sink_wenable;
  reg [32-1:0] _mystream_sum_vec26_sink_wdata;
  reg _mystream_sum_vec26_sink_fifo_enq;
  reg [32-1:0] _mystream_sum_vec26_sink_fifo_wdata;
  reg [32-1:0] _mystream_sum_vec26_sink_immediate;
  reg [33-1:0] _mystream_sum_vec27_sink_count;
  reg [5-1:0] _mystream_sum_vec27_sink_mode;
  reg [16-1:0] _mystream_sum_vec27_sink_generator_id;
  reg [32-1:0] _mystream_sum_vec27_sink_offset;
  reg [33-1:0] _mystream_sum_vec27_sink_size;
  reg [32-1:0] _mystream_sum_vec27_sink_stride;
  reg [32-1:0] _mystream_sum_vec27_sink_offset_buf;
  reg [33-1:0] _mystream_sum_vec27_sink_size_buf;
  reg [32-1:0] _mystream_sum_vec27_sink_stride_buf;
  reg [8-1:0] _mystream_sum_vec27_sink_sel;
  reg [32-1:0] _mystream_sum_vec27_sink_waddr;
  reg _mystream_sum_vec27_sink_wenable;
  reg [32-1:0] _mystream_sum_vec27_sink_wdata;
  reg _mystream_sum_vec27_sink_fifo_enq;
  reg [32-1:0] _mystream_sum_vec27_sink_fifo_wdata;
  reg [32-1:0] _mystream_sum_vec27_sink_immediate;
  reg [33-1:0] _mystream_sum_vec28_sink_count;
  reg [5-1:0] _mystream_sum_vec28_sink_mode;
  reg [16-1:0] _mystream_sum_vec28_sink_generator_id;
  reg [32-1:0] _mystream_sum_vec28_sink_offset;
  reg [33-1:0] _mystream_sum_vec28_sink_size;
  reg [32-1:0] _mystream_sum_vec28_sink_stride;
  reg [32-1:0] _mystream_sum_vec28_sink_offset_buf;
  reg [33-1:0] _mystream_sum_vec28_sink_size_buf;
  reg [32-1:0] _mystream_sum_vec28_sink_stride_buf;
  reg [8-1:0] _mystream_sum_vec28_sink_sel;
  reg [32-1:0] _mystream_sum_vec28_sink_waddr;
  reg _mystream_sum_vec28_sink_wenable;
  reg [32-1:0] _mystream_sum_vec28_sink_wdata;
  reg _mystream_sum_vec28_sink_fifo_enq;
  reg [32-1:0] _mystream_sum_vec28_sink_fifo_wdata;
  reg [32-1:0] _mystream_sum_vec28_sink_immediate;
  reg [33-1:0] _mystream_sum_vec29_sink_count;
  reg [5-1:0] _mystream_sum_vec29_sink_mode;
  reg [16-1:0] _mystream_sum_vec29_sink_generator_id;
  reg [32-1:0] _mystream_sum_vec29_sink_offset;
  reg [33-1:0] _mystream_sum_vec29_sink_size;
  reg [32-1:0] _mystream_sum_vec29_sink_stride;
  reg [32-1:0] _mystream_sum_vec29_sink_offset_buf;
  reg [33-1:0] _mystream_sum_vec29_sink_size_buf;
  reg [32-1:0] _mystream_sum_vec29_sink_stride_buf;
  reg [8-1:0] _mystream_sum_vec29_sink_sel;
  reg [32-1:0] _mystream_sum_vec29_sink_waddr;
  reg _mystream_sum_vec29_sink_wenable;
  reg [32-1:0] _mystream_sum_vec29_sink_wdata;
  reg _mystream_sum_vec29_sink_fifo_enq;
  reg [32-1:0] _mystream_sum_vec29_sink_fifo_wdata;
  reg [32-1:0] _mystream_sum_vec29_sink_immediate;
  reg [33-1:0] _mystream_sum_vec30_sink_count;
  reg [5-1:0] _mystream_sum_vec30_sink_mode;
  reg [16-1:0] _mystream_sum_vec30_sink_generator_id;
  reg [32-1:0] _mystream_sum_vec30_sink_offset;
  reg [33-1:0] _mystream_sum_vec30_sink_size;
  reg [32-1:0] _mystream_sum_vec30_sink_stride;
  reg [32-1:0] _mystream_sum_vec30_sink_offset_buf;
  reg [33-1:0] _mystream_sum_vec30_sink_size_buf;
  reg [32-1:0] _mystream_sum_vec30_sink_stride_buf;
  reg [8-1:0] _mystream_sum_vec30_sink_sel;
  reg [32-1:0] _mystream_sum_vec30_sink_waddr;
  reg _mystream_sum_vec30_sink_wenable;
  reg [32-1:0] _mystream_sum_vec30_sink_wdata;
  reg _mystream_sum_vec30_sink_fifo_enq;
  reg [32-1:0] _mystream_sum_vec30_sink_fifo_wdata;
  reg [32-1:0] _mystream_sum_vec30_sink_immediate;
  reg [33-1:0] _mystream_sum_vec31_sink_count;
  reg [5-1:0] _mystream_sum_vec31_sink_mode;
  reg [16-1:0] _mystream_sum_vec31_sink_generator_id;
  reg [32-1:0] _mystream_sum_vec31_sink_offset;
  reg [33-1:0] _mystream_sum_vec31_sink_size;
  reg [32-1:0] _mystream_sum_vec31_sink_stride;
  reg [32-1:0] _mystream_sum_vec31_sink_offset_buf;
  reg [33-1:0] _mystream_sum_vec31_sink_size_buf;
  reg [32-1:0] _mystream_sum_vec31_sink_stride_buf;
  reg [8-1:0] _mystream_sum_vec31_sink_sel;
  reg [32-1:0] _mystream_sum_vec31_sink_waddr;
  reg _mystream_sum_vec31_sink_wenable;
  reg [32-1:0] _mystream_sum_vec31_sink_wdata;
  reg _mystream_sum_vec31_sink_fifo_enq;
  reg [32-1:0] _mystream_sum_vec31_sink_fifo_wdata;
  reg [32-1:0] _mystream_sum_vec31_sink_immediate;
  reg [32-1:0] counter;
  reg [32-1:0] th_comp;
  localparam th_comp_init = 0;
  reg signed [32-1:0] _th_comp_size_0;
  reg signed [32-1:0] _th_comp_offset_b_1;
  reg signed [32-1:0] _th_comp_offset_2;
  wire [32-1:0] _dma_read_packed_high_local_size_11;
  assign _dma_read_packed_high_local_size_11 = _th_comp_size_0 >> 5;
  wire [5-1:0] _dma_read_packed_low_local_size_12;
  assign _dma_read_packed_low_local_size_12 = _th_comp_size_0 & { 5{ 1'd1 } };
  wire [32-1:0] _dma_read_packed_local_packed_size_13;
  assign _dma_read_packed_local_packed_size_13 = (_dma_read_packed_low_local_size_12 > 0)? _dma_read_packed_high_local_size_11 + 1 : _dma_read_packed_high_local_size_11;
  wire [32-1:0] mask_addr_shifted_14;
  assign mask_addr_shifted_14 = 0 + (_th_comp_size_0 << 2) >> 2;
  wire [32-1:0] mask_addr_masked_15;
  assign mask_addr_masked_15 = mask_addr_shifted_14 << 2;
  reg [32-1:0] _myaxi_read_req_fsm;
  localparam _myaxi_read_req_fsm_init = 0;
  reg [33-1:0] _myaxi_read_cur_global_size;
  reg _myaxi_read_cont;
  wire [8-1:0] pack_read_req_op_sel_16;
  wire [32-1:0] pack_read_req_local_addr_17;
  wire [32-1:0] pack_read_req_local_stride_18;
  wire [33-1:0] pack_read_req_local_size_19;
  wire [32-1:0] pack_read_req_local_blocksize_20;
  assign pack_read_req_op_sel_16 = _myaxi_read_op_sel;
  assign pack_read_req_local_addr_17 = _myaxi_read_local_addr;
  assign pack_read_req_local_stride_18 = _myaxi_read_local_stride;
  assign pack_read_req_local_size_19 = _myaxi_read_local_size;
  assign pack_read_req_local_blocksize_20 = _myaxi_read_local_blocksize;
  wire [137-1:0] pack_read_req_packed_21;
  assign pack_read_req_packed_21 = { pack_read_req_op_sel_16, pack_read_req_local_addr_17, pack_read_req_local_stride_18, pack_read_req_local_size_19, pack_read_req_local_blocksize_20 };
  assign _myaxi_read_req_fifo_wdata = ((_myaxi_read_req_fsm == 0) && _myaxi_read_start && !_myaxi_read_req_fifo_almost_full)? pack_read_req_packed_21 : 'hx;
  assign _myaxi_read_req_fifo_enq = ((_myaxi_read_req_fsm == 0) && _myaxi_read_start && !_myaxi_read_req_fifo_almost_full)? (_myaxi_read_req_fsm == 0) && _myaxi_read_start && !_myaxi_read_req_fifo_almost_full && !_myaxi_read_req_fifo_almost_full : 0;
  localparam _tmp_22 = 1;
  wire [_tmp_22-1:0] _tmp_23;
  assign _tmp_23 = !_myaxi_read_req_fifo_almost_full;
  reg [_tmp_22-1:0] __tmp_23_1;
  wire [32-1:0] mask_addr_shifted_24;
  assign mask_addr_shifted_24 = _myaxi_read_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_25;
  assign mask_addr_masked_25 = mask_addr_shifted_24 << 2;
  wire [32-1:0] mask_addr_shifted_26;
  assign mask_addr_shifted_26 = _myaxi_read_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_27;
  assign mask_addr_masked_27 = mask_addr_shifted_26 << 2;
  wire [32-1:0] mask_addr_shifted_28;
  assign mask_addr_shifted_28 = _myaxi_read_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_29;
  assign mask_addr_masked_29 = mask_addr_shifted_28 << 2;
  wire [32-1:0] mask_addr_shifted_30;
  assign mask_addr_shifted_30 = _myaxi_read_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_31;
  assign mask_addr_masked_31 = mask_addr_shifted_30 << 2;
  wire [32-1:0] mask_addr_shifted_32;
  assign mask_addr_shifted_32 = _myaxi_read_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_33;
  assign mask_addr_masked_33 = mask_addr_shifted_32 << 2;
  wire [32-1:0] mask_addr_shifted_34;
  assign mask_addr_shifted_34 = _myaxi_read_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_35;
  assign mask_addr_masked_35 = mask_addr_shifted_34 << 2;
  reg _myaxi_cond_0_1;
  reg [32-1:0] _myaxi_read_data_narrow_fsm;
  localparam _myaxi_read_data_narrow_fsm_init = 0;
  reg [1024-1:0] _myaxi_read_narrow_wdata_36;
  reg _myaxi_read_narrow_wvalid_37;
  reg [5-1:0] _myaxi_read_narrow_count_38;
  reg [32-1:0] write_burst_packed_fsm_0;
  localparam write_burst_packed_fsm_0_init = 0;
  reg [25-1:0] write_burst_packed_addr_39;
  reg [25-1:0] write_burst_packed_stride_40;
  reg [33-1:0] write_burst_packed_length_41;
  reg write_burst_packed_done_42;
  wire [20-1:0] write_burst_packed_ram_addr_43;
  assign write_burst_packed_ram_addr_43 = write_burst_packed_addr_39 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_44;
  assign write_burst_packed_ram_wdata_44 = _myaxi_read_narrow_wdata_36 >> 0;
  assign ram_a_0_0_wdata = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_wdata_44 : 'hx;
  assign ram_a_0_0_wenable = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_45;
  assign write_burst_packed_ram_addr_45 = write_burst_packed_addr_39 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_46;
  assign write_burst_packed_ram_wdata_46 = _myaxi_read_narrow_wdata_36 >> 32;
  assign ram_a_1_0_wdata = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_wdata_46 : 'hx;
  assign ram_a_1_0_wenable = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_47;
  assign write_burst_packed_ram_addr_47 = write_burst_packed_addr_39 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_48;
  assign write_burst_packed_ram_wdata_48 = _myaxi_read_narrow_wdata_36 >> 64;
  assign ram_a_2_0_wdata = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_wdata_48 : 'hx;
  assign ram_a_2_0_wenable = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_49;
  assign write_burst_packed_ram_addr_49 = write_burst_packed_addr_39 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_50;
  assign write_burst_packed_ram_wdata_50 = _myaxi_read_narrow_wdata_36 >> 96;
  assign ram_a_3_0_wdata = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_wdata_50 : 'hx;
  assign ram_a_3_0_wenable = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_51;
  assign write_burst_packed_ram_addr_51 = write_burst_packed_addr_39 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_52;
  assign write_burst_packed_ram_wdata_52 = _myaxi_read_narrow_wdata_36 >> 128;
  assign ram_a_4_0_wdata = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_wdata_52 : 'hx;
  assign ram_a_4_0_wenable = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_53;
  assign write_burst_packed_ram_addr_53 = write_burst_packed_addr_39 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_54;
  assign write_burst_packed_ram_wdata_54 = _myaxi_read_narrow_wdata_36 >> 160;
  assign ram_a_5_0_wdata = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_wdata_54 : 'hx;
  assign ram_a_5_0_wenable = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_55;
  assign write_burst_packed_ram_addr_55 = write_burst_packed_addr_39 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_56;
  assign write_burst_packed_ram_wdata_56 = _myaxi_read_narrow_wdata_36 >> 192;
  assign ram_a_6_0_wdata = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_wdata_56 : 'hx;
  assign ram_a_6_0_wenable = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_57;
  assign write_burst_packed_ram_addr_57 = write_burst_packed_addr_39 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_58;
  assign write_burst_packed_ram_wdata_58 = _myaxi_read_narrow_wdata_36 >> 224;
  assign ram_a_7_0_wdata = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_wdata_58 : 'hx;
  assign ram_a_7_0_wenable = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_59;
  assign write_burst_packed_ram_addr_59 = write_burst_packed_addr_39 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_60;
  assign write_burst_packed_ram_wdata_60 = _myaxi_read_narrow_wdata_36 >> 256;
  assign ram_a_8_0_wdata = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_wdata_60 : 'hx;
  assign ram_a_8_0_wenable = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_61;
  assign write_burst_packed_ram_addr_61 = write_burst_packed_addr_39 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_62;
  assign write_burst_packed_ram_wdata_62 = _myaxi_read_narrow_wdata_36 >> 288;
  assign ram_a_9_0_wdata = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_wdata_62 : 'hx;
  assign ram_a_9_0_wenable = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_63;
  assign write_burst_packed_ram_addr_63 = write_burst_packed_addr_39 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_64;
  assign write_burst_packed_ram_wdata_64 = _myaxi_read_narrow_wdata_36 >> 320;
  assign ram_a_10_0_wdata = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_wdata_64 : 'hx;
  assign ram_a_10_0_wenable = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_65;
  assign write_burst_packed_ram_addr_65 = write_burst_packed_addr_39 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_66;
  assign write_burst_packed_ram_wdata_66 = _myaxi_read_narrow_wdata_36 >> 352;
  assign ram_a_11_0_wdata = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_wdata_66 : 'hx;
  assign ram_a_11_0_wenable = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_67;
  assign write_burst_packed_ram_addr_67 = write_burst_packed_addr_39 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_68;
  assign write_burst_packed_ram_wdata_68 = _myaxi_read_narrow_wdata_36 >> 384;
  assign ram_a_12_0_wdata = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_wdata_68 : 'hx;
  assign ram_a_12_0_wenable = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_69;
  assign write_burst_packed_ram_addr_69 = write_burst_packed_addr_39 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_70;
  assign write_burst_packed_ram_wdata_70 = _myaxi_read_narrow_wdata_36 >> 416;
  assign ram_a_13_0_wdata = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_wdata_70 : 'hx;
  assign ram_a_13_0_wenable = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_71;
  assign write_burst_packed_ram_addr_71 = write_burst_packed_addr_39 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_72;
  assign write_burst_packed_ram_wdata_72 = _myaxi_read_narrow_wdata_36 >> 448;
  assign ram_a_14_0_wdata = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_wdata_72 : 'hx;
  assign ram_a_14_0_wenable = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_73;
  assign write_burst_packed_ram_addr_73 = write_burst_packed_addr_39 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_74;
  assign write_burst_packed_ram_wdata_74 = _myaxi_read_narrow_wdata_36 >> 480;
  assign ram_a_15_0_wdata = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_wdata_74 : 'hx;
  assign ram_a_15_0_wenable = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_75;
  assign write_burst_packed_ram_addr_75 = write_burst_packed_addr_39 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_76;
  assign write_burst_packed_ram_wdata_76 = _myaxi_read_narrow_wdata_36 >> 512;
  assign ram_a_16_0_wdata = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_wdata_76 : 'hx;
  assign ram_a_16_0_wenable = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_77;
  assign write_burst_packed_ram_addr_77 = write_burst_packed_addr_39 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_78;
  assign write_burst_packed_ram_wdata_78 = _myaxi_read_narrow_wdata_36 >> 544;
  assign ram_a_17_0_wdata = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_wdata_78 : 'hx;
  assign ram_a_17_0_wenable = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_79;
  assign write_burst_packed_ram_addr_79 = write_burst_packed_addr_39 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_80;
  assign write_burst_packed_ram_wdata_80 = _myaxi_read_narrow_wdata_36 >> 576;
  assign ram_a_18_0_wdata = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_wdata_80 : 'hx;
  assign ram_a_18_0_wenable = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_81;
  assign write_burst_packed_ram_addr_81 = write_burst_packed_addr_39 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_82;
  assign write_burst_packed_ram_wdata_82 = _myaxi_read_narrow_wdata_36 >> 608;
  assign ram_a_19_0_wdata = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_wdata_82 : 'hx;
  assign ram_a_19_0_wenable = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_83;
  assign write_burst_packed_ram_addr_83 = write_burst_packed_addr_39 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_84;
  assign write_burst_packed_ram_wdata_84 = _myaxi_read_narrow_wdata_36 >> 640;
  assign ram_a_20_0_wdata = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_wdata_84 : 'hx;
  assign ram_a_20_0_wenable = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_85;
  assign write_burst_packed_ram_addr_85 = write_burst_packed_addr_39 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_86;
  assign write_burst_packed_ram_wdata_86 = _myaxi_read_narrow_wdata_36 >> 672;
  assign ram_a_21_0_wdata = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_wdata_86 : 'hx;
  assign ram_a_21_0_wenable = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_87;
  assign write_burst_packed_ram_addr_87 = write_burst_packed_addr_39 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_88;
  assign write_burst_packed_ram_wdata_88 = _myaxi_read_narrow_wdata_36 >> 704;
  assign ram_a_22_0_wdata = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_wdata_88 : 'hx;
  assign ram_a_22_0_wenable = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_89;
  assign write_burst_packed_ram_addr_89 = write_burst_packed_addr_39 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_90;
  assign write_burst_packed_ram_wdata_90 = _myaxi_read_narrow_wdata_36 >> 736;
  assign ram_a_23_0_wdata = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_wdata_90 : 'hx;
  assign ram_a_23_0_wenable = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_91;
  assign write_burst_packed_ram_addr_91 = write_burst_packed_addr_39 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_92;
  assign write_burst_packed_ram_wdata_92 = _myaxi_read_narrow_wdata_36 >> 768;
  assign ram_a_24_0_wdata = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_wdata_92 : 'hx;
  assign ram_a_24_0_wenable = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_93;
  assign write_burst_packed_ram_addr_93 = write_burst_packed_addr_39 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_94;
  assign write_burst_packed_ram_wdata_94 = _myaxi_read_narrow_wdata_36 >> 800;
  assign ram_a_25_0_wdata = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_wdata_94 : 'hx;
  assign ram_a_25_0_wenable = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_95;
  assign write_burst_packed_ram_addr_95 = write_burst_packed_addr_39 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_96;
  assign write_burst_packed_ram_wdata_96 = _myaxi_read_narrow_wdata_36 >> 832;
  assign ram_a_26_0_wdata = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_wdata_96 : 'hx;
  assign ram_a_26_0_wenable = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_97;
  assign write_burst_packed_ram_addr_97 = write_burst_packed_addr_39 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_98;
  assign write_burst_packed_ram_wdata_98 = _myaxi_read_narrow_wdata_36 >> 864;
  assign ram_a_27_0_wdata = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_wdata_98 : 'hx;
  assign ram_a_27_0_wenable = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_99;
  assign write_burst_packed_ram_addr_99 = write_burst_packed_addr_39 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_100;
  assign write_burst_packed_ram_wdata_100 = _myaxi_read_narrow_wdata_36 >> 896;
  assign ram_a_28_0_wdata = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_wdata_100 : 'hx;
  assign ram_a_28_0_wenable = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_101;
  assign write_burst_packed_ram_addr_101 = write_burst_packed_addr_39 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_102;
  assign write_burst_packed_ram_wdata_102 = _myaxi_read_narrow_wdata_36 >> 928;
  assign ram_a_29_0_wdata = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_wdata_102 : 'hx;
  assign ram_a_29_0_wenable = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_103;
  assign write_burst_packed_ram_addr_103 = write_burst_packed_addr_39 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_104;
  assign write_burst_packed_ram_wdata_104 = _myaxi_read_narrow_wdata_36 >> 960;
  assign ram_a_30_0_wdata = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_wdata_104 : 'hx;
  assign ram_a_30_0_wenable = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_105;
  assign write_burst_packed_ram_addr_105 = write_burst_packed_addr_39 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_106;
  assign write_burst_packed_ram_wdata_106 = _myaxi_read_narrow_wdata_36 >> 992;
  assign ram_a_31_0_wdata = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_wdata_106 : 'hx;
  assign ram_a_31_0_wenable = ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  wire [32-1:0] _dma_read_packed_high_local_size_107;
  assign _dma_read_packed_high_local_size_107 = _th_comp_size_0 >> 5;
  wire [5-1:0] _dma_read_packed_low_local_size_108;
  assign _dma_read_packed_low_local_size_108 = _th_comp_size_0 & { 5{ 1'd1 } };
  wire [32-1:0] _dma_read_packed_local_packed_size_109;
  assign _dma_read_packed_local_packed_size_109 = (_dma_read_packed_low_local_size_108 > 0)? _dma_read_packed_high_local_size_107 + 1 : _dma_read_packed_high_local_size_107;
  wire [32-1:0] mask_addr_shifted_110;
  assign mask_addr_shifted_110 = _th_comp_offset_b_1 + (_th_comp_size_0 << 2) >> 2;
  wire [32-1:0] mask_addr_masked_111;
  assign mask_addr_masked_111 = mask_addr_shifted_110 << 2;
  reg [1024-1:0] _myaxi_read_narrow_wdata_112;
  reg _myaxi_read_narrow_wvalid_113;
  reg [5-1:0] _myaxi_read_narrow_count_114;
  reg [32-1:0] write_burst_packed_fsm_1;
  localparam write_burst_packed_fsm_1_init = 0;
  reg [25-1:0] write_burst_packed_addr_115;
  reg [25-1:0] write_burst_packed_stride_116;
  reg [33-1:0] write_burst_packed_length_117;
  reg write_burst_packed_done_118;
  wire [20-1:0] write_burst_packed_ram_addr_119;
  assign write_burst_packed_ram_addr_119 = write_burst_packed_addr_115 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_120;
  assign write_burst_packed_ram_wdata_120 = _myaxi_read_narrow_wdata_112 >> 0;
  assign ram_b_0_0_wdata = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_wdata_120 : 'hx;
  assign ram_b_0_0_wenable = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_121;
  assign write_burst_packed_ram_addr_121 = write_burst_packed_addr_115 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_122;
  assign write_burst_packed_ram_wdata_122 = _myaxi_read_narrow_wdata_112 >> 32;
  assign ram_b_1_0_wdata = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_wdata_122 : 'hx;
  assign ram_b_1_0_wenable = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_123;
  assign write_burst_packed_ram_addr_123 = write_burst_packed_addr_115 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_124;
  assign write_burst_packed_ram_wdata_124 = _myaxi_read_narrow_wdata_112 >> 64;
  assign ram_b_2_0_wdata = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_wdata_124 : 'hx;
  assign ram_b_2_0_wenable = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_125;
  assign write_burst_packed_ram_addr_125 = write_burst_packed_addr_115 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_126;
  assign write_burst_packed_ram_wdata_126 = _myaxi_read_narrow_wdata_112 >> 96;
  assign ram_b_3_0_wdata = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_wdata_126 : 'hx;
  assign ram_b_3_0_wenable = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_127;
  assign write_burst_packed_ram_addr_127 = write_burst_packed_addr_115 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_128;
  assign write_burst_packed_ram_wdata_128 = _myaxi_read_narrow_wdata_112 >> 128;
  assign ram_b_4_0_wdata = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_wdata_128 : 'hx;
  assign ram_b_4_0_wenable = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_129;
  assign write_burst_packed_ram_addr_129 = write_burst_packed_addr_115 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_130;
  assign write_burst_packed_ram_wdata_130 = _myaxi_read_narrow_wdata_112 >> 160;
  assign ram_b_5_0_wdata = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_wdata_130 : 'hx;
  assign ram_b_5_0_wenable = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_131;
  assign write_burst_packed_ram_addr_131 = write_burst_packed_addr_115 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_132;
  assign write_burst_packed_ram_wdata_132 = _myaxi_read_narrow_wdata_112 >> 192;
  assign ram_b_6_0_wdata = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_wdata_132 : 'hx;
  assign ram_b_6_0_wenable = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_133;
  assign write_burst_packed_ram_addr_133 = write_burst_packed_addr_115 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_134;
  assign write_burst_packed_ram_wdata_134 = _myaxi_read_narrow_wdata_112 >> 224;
  assign ram_b_7_0_wdata = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_wdata_134 : 'hx;
  assign ram_b_7_0_wenable = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_135;
  assign write_burst_packed_ram_addr_135 = write_burst_packed_addr_115 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_136;
  assign write_burst_packed_ram_wdata_136 = _myaxi_read_narrow_wdata_112 >> 256;
  assign ram_b_8_0_wdata = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_wdata_136 : 'hx;
  assign ram_b_8_0_wenable = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_137;
  assign write_burst_packed_ram_addr_137 = write_burst_packed_addr_115 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_138;
  assign write_burst_packed_ram_wdata_138 = _myaxi_read_narrow_wdata_112 >> 288;
  assign ram_b_9_0_wdata = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_wdata_138 : 'hx;
  assign ram_b_9_0_wenable = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_139;
  assign write_burst_packed_ram_addr_139 = write_burst_packed_addr_115 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_140;
  assign write_burst_packed_ram_wdata_140 = _myaxi_read_narrow_wdata_112 >> 320;
  assign ram_b_10_0_wdata = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_wdata_140 : 'hx;
  assign ram_b_10_0_wenable = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_141;
  assign write_burst_packed_ram_addr_141 = write_burst_packed_addr_115 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_142;
  assign write_burst_packed_ram_wdata_142 = _myaxi_read_narrow_wdata_112 >> 352;
  assign ram_b_11_0_wdata = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_wdata_142 : 'hx;
  assign ram_b_11_0_wenable = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_143;
  assign write_burst_packed_ram_addr_143 = write_burst_packed_addr_115 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_144;
  assign write_burst_packed_ram_wdata_144 = _myaxi_read_narrow_wdata_112 >> 384;
  assign ram_b_12_0_wdata = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_wdata_144 : 'hx;
  assign ram_b_12_0_wenable = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_145;
  assign write_burst_packed_ram_addr_145 = write_burst_packed_addr_115 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_146;
  assign write_burst_packed_ram_wdata_146 = _myaxi_read_narrow_wdata_112 >> 416;
  assign ram_b_13_0_wdata = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_wdata_146 : 'hx;
  assign ram_b_13_0_wenable = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_147;
  assign write_burst_packed_ram_addr_147 = write_burst_packed_addr_115 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_148;
  assign write_burst_packed_ram_wdata_148 = _myaxi_read_narrow_wdata_112 >> 448;
  assign ram_b_14_0_wdata = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_wdata_148 : 'hx;
  assign ram_b_14_0_wenable = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_149;
  assign write_burst_packed_ram_addr_149 = write_burst_packed_addr_115 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_150;
  assign write_burst_packed_ram_wdata_150 = _myaxi_read_narrow_wdata_112 >> 480;
  assign ram_b_15_0_wdata = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_wdata_150 : 'hx;
  assign ram_b_15_0_wenable = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_151;
  assign write_burst_packed_ram_addr_151 = write_burst_packed_addr_115 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_152;
  assign write_burst_packed_ram_wdata_152 = _myaxi_read_narrow_wdata_112 >> 512;
  assign ram_b_16_0_wdata = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_wdata_152 : 'hx;
  assign ram_b_16_0_wenable = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_153;
  assign write_burst_packed_ram_addr_153 = write_burst_packed_addr_115 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_154;
  assign write_burst_packed_ram_wdata_154 = _myaxi_read_narrow_wdata_112 >> 544;
  assign ram_b_17_0_wdata = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_wdata_154 : 'hx;
  assign ram_b_17_0_wenable = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_155;
  assign write_burst_packed_ram_addr_155 = write_burst_packed_addr_115 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_156;
  assign write_burst_packed_ram_wdata_156 = _myaxi_read_narrow_wdata_112 >> 576;
  assign ram_b_18_0_wdata = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_wdata_156 : 'hx;
  assign ram_b_18_0_wenable = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_157;
  assign write_burst_packed_ram_addr_157 = write_burst_packed_addr_115 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_158;
  assign write_burst_packed_ram_wdata_158 = _myaxi_read_narrow_wdata_112 >> 608;
  assign ram_b_19_0_wdata = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_wdata_158 : 'hx;
  assign ram_b_19_0_wenable = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_159;
  assign write_burst_packed_ram_addr_159 = write_burst_packed_addr_115 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_160;
  assign write_burst_packed_ram_wdata_160 = _myaxi_read_narrow_wdata_112 >> 640;
  assign ram_b_20_0_wdata = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_wdata_160 : 'hx;
  assign ram_b_20_0_wenable = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_161;
  assign write_burst_packed_ram_addr_161 = write_burst_packed_addr_115 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_162;
  assign write_burst_packed_ram_wdata_162 = _myaxi_read_narrow_wdata_112 >> 672;
  assign ram_b_21_0_wdata = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_wdata_162 : 'hx;
  assign ram_b_21_0_wenable = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_163;
  assign write_burst_packed_ram_addr_163 = write_burst_packed_addr_115 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_164;
  assign write_burst_packed_ram_wdata_164 = _myaxi_read_narrow_wdata_112 >> 704;
  assign ram_b_22_0_wdata = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_wdata_164 : 'hx;
  assign ram_b_22_0_wenable = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_165;
  assign write_burst_packed_ram_addr_165 = write_burst_packed_addr_115 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_166;
  assign write_burst_packed_ram_wdata_166 = _myaxi_read_narrow_wdata_112 >> 736;
  assign ram_b_23_0_wdata = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_wdata_166 : 'hx;
  assign ram_b_23_0_wenable = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_167;
  assign write_burst_packed_ram_addr_167 = write_burst_packed_addr_115 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_168;
  assign write_burst_packed_ram_wdata_168 = _myaxi_read_narrow_wdata_112 >> 768;
  assign ram_b_24_0_wdata = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_wdata_168 : 'hx;
  assign ram_b_24_0_wenable = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_169;
  assign write_burst_packed_ram_addr_169 = write_burst_packed_addr_115 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_170;
  assign write_burst_packed_ram_wdata_170 = _myaxi_read_narrow_wdata_112 >> 800;
  assign ram_b_25_0_wdata = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_wdata_170 : 'hx;
  assign ram_b_25_0_wenable = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_171;
  assign write_burst_packed_ram_addr_171 = write_burst_packed_addr_115 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_172;
  assign write_burst_packed_ram_wdata_172 = _myaxi_read_narrow_wdata_112 >> 832;
  assign ram_b_26_0_wdata = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_wdata_172 : 'hx;
  assign ram_b_26_0_wenable = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_173;
  assign write_burst_packed_ram_addr_173 = write_burst_packed_addr_115 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_174;
  assign write_burst_packed_ram_wdata_174 = _myaxi_read_narrow_wdata_112 >> 864;
  assign ram_b_27_0_wdata = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_wdata_174 : 'hx;
  assign ram_b_27_0_wenable = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_175;
  assign write_burst_packed_ram_addr_175 = write_burst_packed_addr_115 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_176;
  assign write_burst_packed_ram_wdata_176 = _myaxi_read_narrow_wdata_112 >> 896;
  assign ram_b_28_0_wdata = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_wdata_176 : 'hx;
  assign ram_b_28_0_wenable = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_177;
  assign write_burst_packed_ram_addr_177 = write_burst_packed_addr_115 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_178;
  assign write_burst_packed_ram_wdata_178 = _myaxi_read_narrow_wdata_112 >> 928;
  assign ram_b_29_0_wdata = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_wdata_178 : 'hx;
  assign ram_b_29_0_wenable = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_179;
  assign write_burst_packed_ram_addr_179 = write_burst_packed_addr_115 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_180;
  assign write_burst_packed_ram_wdata_180 = _myaxi_read_narrow_wdata_112 >> 960;
  assign ram_b_30_0_wdata = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_wdata_180 : 'hx;
  assign ram_b_30_0_wenable = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_181;
  assign write_burst_packed_ram_addr_181 = write_burst_packed_addr_115 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_182;
  assign write_burst_packed_ram_wdata_182 = _myaxi_read_narrow_wdata_112 >> 992;
  assign ram_b_31_0_wdata = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_wdata_182 : 'hx;
  assign ram_b_31_0_wenable = ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  reg signed [32-1:0] _th_comp_size_3;
  reg signed [32-1:0] _th_comp_offset_4;
  reg signed [32-1:0] _th_comp_start_time_5;
  wire signed [32-1:0] mystream_size_data;
  wire signed [32-1:0] mystream_tensor_size_data;
  wire signed [32-1:0] mystream_a0_data;
  wire signed [32-1:0] mystream_a1_data;
  wire signed [32-1:0] mystream_a2_data;
  wire signed [32-1:0] mystream_a3_data;
  wire signed [32-1:0] mystream_a4_data;
  wire signed [32-1:0] mystream_a5_data;
  wire signed [32-1:0] mystream_a6_data;
  wire signed [32-1:0] mystream_a7_data;
  wire signed [32-1:0] mystream_a8_data;
  wire signed [32-1:0] mystream_a9_data;
  wire signed [32-1:0] mystream_a10_data;
  wire signed [32-1:0] mystream_a11_data;
  wire signed [32-1:0] mystream_a12_data;
  wire signed [32-1:0] mystream_a13_data;
  wire signed [32-1:0] mystream_a14_data;
  wire signed [32-1:0] mystream_a15_data;
  wire signed [32-1:0] mystream_a16_data;
  wire signed [32-1:0] mystream_a17_data;
  wire signed [32-1:0] mystream_a18_data;
  wire signed [32-1:0] mystream_a19_data;
  wire signed [32-1:0] mystream_a20_data;
  wire signed [32-1:0] mystream_a21_data;
  wire signed [32-1:0] mystream_a22_data;
  wire signed [32-1:0] mystream_a23_data;
  wire signed [32-1:0] mystream_a24_data;
  wire signed [32-1:0] mystream_a25_data;
  wire signed [32-1:0] mystream_a26_data;
  wire signed [32-1:0] mystream_a27_data;
  wire signed [32-1:0] mystream_a28_data;
  wire signed [32-1:0] mystream_a29_data;
  wire signed [32-1:0] mystream_a30_data;
  wire signed [32-1:0] mystream_a31_data;
  wire signed [32-1:0] mystream_b0_data;
  wire signed [32-1:0] mystream_b1_data;
  wire signed [32-1:0] mystream_b2_data;
  wire signed [32-1:0] mystream_b3_data;
  wire signed [32-1:0] mystream_b4_data;
  wire signed [32-1:0] mystream_b5_data;
  wire signed [32-1:0] mystream_b6_data;
  wire signed [32-1:0] mystream_b7_data;
  wire signed [32-1:0] mystream_b8_data;
  wire signed [32-1:0] mystream_b9_data;
  wire signed [32-1:0] mystream_b10_data;
  wire signed [32-1:0] mystream_b11_data;
  wire signed [32-1:0] mystream_b12_data;
  wire signed [32-1:0] mystream_b13_data;
  wire signed [32-1:0] mystream_b14_data;
  wire signed [32-1:0] mystream_b15_data;
  wire signed [32-1:0] mystream_b16_data;
  wire signed [32-1:0] mystream_b17_data;
  wire signed [32-1:0] mystream_b18_data;
  wire signed [32-1:0] mystream_b19_data;
  wire signed [32-1:0] mystream_b20_data;
  wire signed [32-1:0] mystream_b21_data;
  wire signed [32-1:0] mystream_b22_data;
  wire signed [32-1:0] mystream_b23_data;
  wire signed [32-1:0] mystream_b24_data;
  wire signed [32-1:0] mystream_b25_data;
  wire signed [32-1:0] mystream_b26_data;
  wire signed [32-1:0] mystream_b27_data;
  wire signed [32-1:0] mystream_b28_data;
  wire signed [32-1:0] mystream_b29_data;
  wire signed [32-1:0] mystream_b30_data;
  wire signed [32-1:0] mystream_b31_data;
  wire signed [32-1:0] mystream_bias0_data;
  wire signed [32-1:0] mystream_bias1_data;
  wire signed [32-1:0] mystream_bias2_data;
  wire signed [32-1:0] mystream_bias3_data;
  wire signed [32-1:0] mystream_bias4_data;
  wire signed [32-1:0] mystream_bias5_data;
  wire signed [32-1:0] mystream_bias6_data;
  wire signed [32-1:0] mystream_bias7_data;
  wire signed [32-1:0] mystream_bias8_data;
  wire signed [32-1:0] mystream_bias9_data;
  wire signed [32-1:0] mystream_bias10_data;
  wire signed [32-1:0] mystream_bias11_data;
  wire signed [32-1:0] mystream_bias12_data;
  wire signed [32-1:0] mystream_bias13_data;
  wire signed [32-1:0] mystream_bias14_data;
  wire signed [32-1:0] mystream_bias15_data;
  wire signed [32-1:0] mystream_bias16_data;
  wire signed [32-1:0] mystream_bias17_data;
  wire signed [32-1:0] mystream_bias18_data;
  wire signed [32-1:0] mystream_bias19_data;
  wire signed [32-1:0] mystream_bias20_data;
  wire signed [32-1:0] mystream_bias21_data;
  wire signed [32-1:0] mystream_bias22_data;
  wire signed [32-1:0] mystream_bias23_data;
  wire signed [32-1:0] mystream_bias24_data;
  wire signed [32-1:0] mystream_bias25_data;
  wire signed [32-1:0] mystream_bias26_data;
  wire signed [32-1:0] mystream_bias27_data;
  wire signed [32-1:0] mystream_bias28_data;
  wire signed [32-1:0] mystream_bias29_data;
  wire signed [32-1:0] mystream_bias30_data;
  wire signed [32-1:0] mystream_bias31_data;
  wire [1-1:0] mystream__reduce_reset_data;
  reg __mystream_stream_ivalid_1;
  reg __mystream_stream_ivalid_2;
  reg __mystream_stream_ivalid_3;
  reg __mystream_stream_ivalid_4;
  reg signed [32-1:0] _plus_data_98;
  reg signed [32-1:0] _plus_data_99;
  reg signed [32-1:0] _plus_data_100;
  reg signed [32-1:0] _plus_data_101;
  reg signed [32-1:0] _plus_data_102;
  reg signed [32-1:0] _plus_data_103;
  reg signed [32-1:0] _plus_data_104;
  reg signed [32-1:0] _plus_data_105;
  reg signed [32-1:0] _plus_data_106;
  reg signed [32-1:0] _plus_data_107;
  reg signed [32-1:0] _plus_data_108;
  reg signed [32-1:0] _plus_data_109;
  reg signed [32-1:0] _plus_data_110;
  reg signed [32-1:0] _plus_data_111;
  reg signed [32-1:0] _plus_data_112;
  reg signed [32-1:0] _plus_data_113;
  reg signed [32-1:0] _plus_data_114;
  reg signed [32-1:0] _plus_data_115;
  reg signed [32-1:0] _plus_data_116;
  reg signed [32-1:0] _plus_data_117;
  reg signed [32-1:0] _plus_data_118;
  reg signed [32-1:0] _plus_data_119;
  reg signed [32-1:0] _plus_data_120;
  reg signed [32-1:0] _plus_data_121;
  reg signed [32-1:0] _plus_data_122;
  reg signed [32-1:0] _plus_data_123;
  reg signed [32-1:0] _plus_data_124;
  reg signed [32-1:0] _plus_data_125;
  reg signed [32-1:0] _plus_data_126;
  reg signed [32-1:0] _plus_data_127;
  reg signed [32-1:0] _plus_data_128;
  reg signed [32-1:0] _plus_data_129;
  reg [32-1:0] _counter_data_131;
  reg [32-1:0] _counter_count_131;
  wire _counter_reset_cond_131;
  assign _counter_reset_cond_131 = mystream__reduce_reset_data;
  wire [32-1:0] _counter_current_count_131;
  assign _counter_current_count_131 = (_counter_reset_cond_131)? 1'sd0 : _counter_count_131;
  reg signed [32-1:0] __delay_data_294__variable_1;
  reg [32-1:0] _plus_data_134;
  reg [32-1:0] _plus_data_137;
  reg [32-1:0] _plus_data_140;
  reg [32-1:0] _plus_data_143;
  reg [32-1:0] _plus_data_146;
  reg [32-1:0] _plus_data_149;
  reg [32-1:0] _plus_data_152;
  reg [32-1:0] _plus_data_155;
  reg [32-1:0] _plus_data_158;
  reg [32-1:0] _plus_data_161;
  reg [32-1:0] _plus_data_164;
  reg [32-1:0] _plus_data_167;
  reg [32-1:0] _plus_data_170;
  reg [32-1:0] _plus_data_173;
  reg [32-1:0] _plus_data_176;
  reg [32-1:0] _plus_data_179;
  reg [32-1:0] _plus_data_182;
  reg [32-1:0] _plus_data_185;
  reg [32-1:0] _plus_data_188;
  reg [32-1:0] _plus_data_191;
  reg [32-1:0] _plus_data_194;
  reg [32-1:0] _plus_data_197;
  reg [32-1:0] _plus_data_200;
  reg [32-1:0] _plus_data_203;
  reg [32-1:0] _plus_data_206;
  reg [32-1:0] _plus_data_209;
  reg [32-1:0] _plus_data_212;
  reg [32-1:0] _plus_data_215;
  reg [32-1:0] _plus_data_218;
  reg [32-1:0] _plus_data_221;
  reg [32-1:0] _plus_data_224;
  reg [32-1:0] _plus_data_227;
  reg signed [32-1:0] __delay_data_295__delay_294__variable_1;
  reg signed [32-1:0] __delay_data_296_plus_98;
  reg signed [32-1:0] __delay_data_298_plus_99;
  reg signed [32-1:0] __delay_data_300_plus_100;
  reg signed [32-1:0] __delay_data_302_plus_101;
  reg signed [32-1:0] __delay_data_304_plus_102;
  reg signed [32-1:0] __delay_data_306_plus_103;
  reg signed [32-1:0] __delay_data_308_plus_104;
  reg signed [32-1:0] __delay_data_310_plus_105;
  reg signed [32-1:0] __delay_data_312_plus_106;
  reg signed [32-1:0] __delay_data_314_plus_107;
  reg signed [32-1:0] __delay_data_316_plus_108;
  reg signed [32-1:0] __delay_data_318_plus_109;
  reg signed [32-1:0] __delay_data_320_plus_110;
  reg signed [32-1:0] __delay_data_322_plus_111;
  reg signed [32-1:0] __delay_data_324_plus_112;
  reg signed [32-1:0] __delay_data_326_plus_113;
  reg signed [32-1:0] __delay_data_328_plus_114;
  reg signed [32-1:0] __delay_data_330_plus_115;
  reg signed [32-1:0] __delay_data_332_plus_116;
  reg signed [32-1:0] __delay_data_334_plus_117;
  reg signed [32-1:0] __delay_data_336_plus_118;
  reg signed [32-1:0] __delay_data_338_plus_119;
  reg signed [32-1:0] __delay_data_340_plus_120;
  reg signed [32-1:0] __delay_data_342_plus_121;
  reg signed [32-1:0] __delay_data_344_plus_122;
  reg signed [32-1:0] __delay_data_346_plus_123;
  reg signed [32-1:0] __delay_data_348_plus_124;
  reg signed [32-1:0] __delay_data_350_plus_125;
  reg signed [32-1:0] __delay_data_352_plus_126;
  reg signed [32-1:0] __delay_data_354_plus_127;
  reg signed [32-1:0] __delay_data_356_plus_128;
  reg signed [32-1:0] __delay_data_358_plus_129;
  reg [1-1:0] _greatereq_data_136;
  reg [1-1:0] _greatereq_data_139;
  reg [1-1:0] _greatereq_data_142;
  reg [1-1:0] _greatereq_data_145;
  reg [1-1:0] _greatereq_data_148;
  reg [1-1:0] _greatereq_data_151;
  reg [1-1:0] _greatereq_data_154;
  reg [1-1:0] _greatereq_data_157;
  reg [1-1:0] _greatereq_data_160;
  reg [1-1:0] _greatereq_data_163;
  reg [1-1:0] _greatereq_data_166;
  reg [1-1:0] _greatereq_data_169;
  reg [1-1:0] _greatereq_data_172;
  reg [1-1:0] _greatereq_data_175;
  reg [1-1:0] _greatereq_data_178;
  reg [1-1:0] _greatereq_data_181;
  reg [1-1:0] _greatereq_data_184;
  reg [1-1:0] _greatereq_data_187;
  reg [1-1:0] _greatereq_data_190;
  reg [1-1:0] _greatereq_data_193;
  reg [1-1:0] _greatereq_data_196;
  reg [1-1:0] _greatereq_data_199;
  reg [1-1:0] _greatereq_data_202;
  reg [1-1:0] _greatereq_data_205;
  reg [1-1:0] _greatereq_data_208;
  reg [1-1:0] _greatereq_data_211;
  reg [1-1:0] _greatereq_data_214;
  reg [1-1:0] _greatereq_data_217;
  reg [1-1:0] _greatereq_data_220;
  reg [1-1:0] _greatereq_data_223;
  reg [1-1:0] _greatereq_data_226;
  reg [1-1:0] _greatereq_data_229;
  reg signed [32-1:0] __delay_data_297__delay_296_plus_98;
  reg signed [32-1:0] __delay_data_299__delay_298_plus_99;
  reg signed [32-1:0] __delay_data_301__delay_300_plus_100;
  reg signed [32-1:0] __delay_data_303__delay_302_plus_101;
  reg signed [32-1:0] __delay_data_305__delay_304_plus_102;
  reg signed [32-1:0] __delay_data_307__delay_306_plus_103;
  reg signed [32-1:0] __delay_data_309__delay_308_plus_104;
  reg signed [32-1:0] __delay_data_311__delay_310_plus_105;
  reg signed [32-1:0] __delay_data_313__delay_312_plus_106;
  reg signed [32-1:0] __delay_data_315__delay_314_plus_107;
  reg signed [32-1:0] __delay_data_317__delay_316_plus_108;
  reg signed [32-1:0] __delay_data_319__delay_318_plus_109;
  reg signed [32-1:0] __delay_data_321__delay_320_plus_110;
  reg signed [32-1:0] __delay_data_323__delay_322_plus_111;
  reg signed [32-1:0] __delay_data_325__delay_324_plus_112;
  reg signed [32-1:0] __delay_data_327__delay_326_plus_113;
  reg signed [32-1:0] __delay_data_329__delay_328_plus_114;
  reg signed [32-1:0] __delay_data_331__delay_330_plus_115;
  reg signed [32-1:0] __delay_data_333__delay_332_plus_116;
  reg signed [32-1:0] __delay_data_335__delay_334_plus_117;
  reg signed [32-1:0] __delay_data_337__delay_336_plus_118;
  reg signed [32-1:0] __delay_data_339__delay_338_plus_119;
  reg signed [32-1:0] __delay_data_341__delay_340_plus_120;
  reg signed [32-1:0] __delay_data_343__delay_342_plus_121;
  reg signed [32-1:0] __delay_data_345__delay_344_plus_122;
  reg signed [32-1:0] __delay_data_347__delay_346_plus_123;
  reg signed [32-1:0] __delay_data_349__delay_348_plus_124;
  reg signed [32-1:0] __delay_data_351__delay_350_plus_125;
  reg signed [32-1:0] __delay_data_353__delay_352_plus_126;
  reg signed [32-1:0] __delay_data_355__delay_354_plus_127;
  reg signed [32-1:0] __delay_data_357__delay_356_plus_128;
  reg signed [32-1:0] __delay_data_359__delay_358_plus_129;
  reg signed [32-1:0] _cond_data_230;
  reg signed [32-1:0] _cond_data_232;
  reg signed [32-1:0] _cond_data_234;
  reg signed [32-1:0] _cond_data_236;
  reg signed [32-1:0] _cond_data_238;
  reg signed [32-1:0] _cond_data_240;
  reg signed [32-1:0] _cond_data_242;
  reg signed [32-1:0] _cond_data_244;
  reg signed [32-1:0] _cond_data_246;
  reg signed [32-1:0] _cond_data_248;
  reg signed [32-1:0] _cond_data_250;
  reg signed [32-1:0] _cond_data_252;
  reg signed [32-1:0] _cond_data_254;
  reg signed [32-1:0] _cond_data_256;
  reg signed [32-1:0] _cond_data_258;
  reg signed [32-1:0] _cond_data_260;
  reg signed [32-1:0] _cond_data_262;
  reg signed [32-1:0] _cond_data_264;
  reg signed [32-1:0] _cond_data_266;
  reg signed [32-1:0] _cond_data_268;
  reg signed [32-1:0] _cond_data_270;
  reg signed [32-1:0] _cond_data_272;
  reg signed [32-1:0] _cond_data_274;
  reg signed [32-1:0] _cond_data_276;
  reg signed [32-1:0] _cond_data_278;
  reg signed [32-1:0] _cond_data_280;
  reg signed [32-1:0] _cond_data_282;
  reg signed [32-1:0] _cond_data_284;
  reg signed [32-1:0] _cond_data_286;
  reg signed [32-1:0] _cond_data_288;
  reg signed [32-1:0] _cond_data_290;
  reg signed [32-1:0] _cond_data_292;
  wire signed [32-1:0] mystream_sum_vec0_data;
  assign mystream_sum_vec0_data = _cond_data_230;
  wire signed [32-1:0] mystream_sum_vec1_data;
  assign mystream_sum_vec1_data = _cond_data_232;
  wire signed [32-1:0] mystream_sum_vec2_data;
  assign mystream_sum_vec2_data = _cond_data_234;
  wire signed [32-1:0] mystream_sum_vec3_data;
  assign mystream_sum_vec3_data = _cond_data_236;
  wire signed [32-1:0] mystream_sum_vec4_data;
  assign mystream_sum_vec4_data = _cond_data_238;
  wire signed [32-1:0] mystream_sum_vec5_data;
  assign mystream_sum_vec5_data = _cond_data_240;
  wire signed [32-1:0] mystream_sum_vec6_data;
  assign mystream_sum_vec6_data = _cond_data_242;
  wire signed [32-1:0] mystream_sum_vec7_data;
  assign mystream_sum_vec7_data = _cond_data_244;
  wire signed [32-1:0] mystream_sum_vec8_data;
  assign mystream_sum_vec8_data = _cond_data_246;
  wire signed [32-1:0] mystream_sum_vec9_data;
  assign mystream_sum_vec9_data = _cond_data_248;
  wire signed [32-1:0] mystream_sum_vec10_data;
  assign mystream_sum_vec10_data = _cond_data_250;
  wire signed [32-1:0] mystream_sum_vec11_data;
  assign mystream_sum_vec11_data = _cond_data_252;
  wire signed [32-1:0] mystream_sum_vec12_data;
  assign mystream_sum_vec12_data = _cond_data_254;
  wire signed [32-1:0] mystream_sum_vec13_data;
  assign mystream_sum_vec13_data = _cond_data_256;
  wire signed [32-1:0] mystream_sum_vec14_data;
  assign mystream_sum_vec14_data = _cond_data_258;
  wire signed [32-1:0] mystream_sum_vec15_data;
  assign mystream_sum_vec15_data = _cond_data_260;
  wire signed [32-1:0] mystream_sum_vec16_data;
  assign mystream_sum_vec16_data = _cond_data_262;
  wire signed [32-1:0] mystream_sum_vec17_data;
  assign mystream_sum_vec17_data = _cond_data_264;
  wire signed [32-1:0] mystream_sum_vec18_data;
  assign mystream_sum_vec18_data = _cond_data_266;
  wire signed [32-1:0] mystream_sum_vec19_data;
  assign mystream_sum_vec19_data = _cond_data_268;
  wire signed [32-1:0] mystream_sum_vec20_data;
  assign mystream_sum_vec20_data = _cond_data_270;
  wire signed [32-1:0] mystream_sum_vec21_data;
  assign mystream_sum_vec21_data = _cond_data_272;
  wire signed [32-1:0] mystream_sum_vec22_data;
  assign mystream_sum_vec22_data = _cond_data_274;
  wire signed [32-1:0] mystream_sum_vec23_data;
  assign mystream_sum_vec23_data = _cond_data_276;
  wire signed [32-1:0] mystream_sum_vec24_data;
  assign mystream_sum_vec24_data = _cond_data_278;
  wire signed [32-1:0] mystream_sum_vec25_data;
  assign mystream_sum_vec25_data = _cond_data_280;
  wire signed [32-1:0] mystream_sum_vec26_data;
  assign mystream_sum_vec26_data = _cond_data_282;
  wire signed [32-1:0] mystream_sum_vec27_data;
  assign mystream_sum_vec27_data = _cond_data_284;
  wire signed [32-1:0] mystream_sum_vec28_data;
  assign mystream_sum_vec28_data = _cond_data_286;
  wire signed [32-1:0] mystream_sum_vec29_data;
  assign mystream_sum_vec29_data = _cond_data_288;
  wire signed [32-1:0] mystream_sum_vec30_data;
  assign mystream_sum_vec30_data = _cond_data_290;
  wire signed [32-1:0] mystream_sum_vec31_data;
  assign mystream_sum_vec31_data = _cond_data_292;
  wire _set_flag_183;
  assign _set_flag_183 = th_comp == 10;
  reg signed [32-1:0] __variable_wdata_1;
  assign mystream_tensor_size_data = __variable_wdata_1;
  wire _set_flag_184;
  assign _set_flag_184 = th_comp == 11;
  reg signed [32-1:0] __variable_wdata_0;
  assign mystream_size_data = __variable_wdata_0;
  reg signed [32-1:0] _th_comp_end_time_6;
  wire _set_flag_185;
  assign _set_flag_185 = th_comp == 14;
  assign ram_a_0_0_addr = (_mystream_stream_oready && _mystream_a0_source_ram_renable && (_mystream_a0_source_sel == 1))? _mystream_a0_source_ram_raddr : 
                          ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_addr_43 : 'hx;
  assign ram_a_0_0_enable = (_mystream_stream_oready && _mystream_a0_source_ram_renable && (_mystream_a0_source_sel == 1))? 1'd1 : 
                            ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  localparam _tmp_186 = 1;
  wire [_tmp_186-1:0] _tmp_187;
  assign _tmp_187 = _mystream_stream_oready && _mystream_a0_source_ram_renable && (_mystream_a0_source_sel == 1);
  reg [_tmp_186-1:0] __tmp_187_1;
  assign _mystream_a0_source_ram_rdata = (_mystream_a0_source_sel == 1)? ram_a_0_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_2;
  assign mystream_a0_data = __variable_wdata_2;
  reg [32-1:0] _mystream_a0_source_fsm_0;
  localparam _mystream_a0_source_fsm_0_init = 0;
  wire _set_flag_188;
  assign _set_flag_188 = th_comp == 15;
  assign ram_a_1_0_addr = (_mystream_stream_oready && _mystream_a1_source_ram_renable && (_mystream_a1_source_sel == 2))? _mystream_a1_source_ram_raddr : 
                          ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_addr_45 : 'hx;
  assign ram_a_1_0_enable = (_mystream_stream_oready && _mystream_a1_source_ram_renable && (_mystream_a1_source_sel == 2))? 1'd1 : 
                            ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  localparam _tmp_189 = 1;
  wire [_tmp_189-1:0] _tmp_190;
  assign _tmp_190 = _mystream_stream_oready && _mystream_a1_source_ram_renable && (_mystream_a1_source_sel == 2);
  reg [_tmp_189-1:0] __tmp_190_1;
  assign _mystream_a1_source_ram_rdata = (_mystream_a1_source_sel == 2)? ram_a_1_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_3;
  assign mystream_a1_data = __variable_wdata_3;
  reg [32-1:0] _mystream_a1_source_fsm_1;
  localparam _mystream_a1_source_fsm_1_init = 0;
  wire _set_flag_191;
  assign _set_flag_191 = th_comp == 16;
  assign ram_a_2_0_addr = (_mystream_stream_oready && _mystream_a2_source_ram_renable && (_mystream_a2_source_sel == 3))? _mystream_a2_source_ram_raddr : 
                          ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_addr_47 : 'hx;
  assign ram_a_2_0_enable = (_mystream_stream_oready && _mystream_a2_source_ram_renable && (_mystream_a2_source_sel == 3))? 1'd1 : 
                            ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  localparam _tmp_192 = 1;
  wire [_tmp_192-1:0] _tmp_193;
  assign _tmp_193 = _mystream_stream_oready && _mystream_a2_source_ram_renable && (_mystream_a2_source_sel == 3);
  reg [_tmp_192-1:0] __tmp_193_1;
  assign _mystream_a2_source_ram_rdata = (_mystream_a2_source_sel == 3)? ram_a_2_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_4;
  assign mystream_a2_data = __variable_wdata_4;
  reg [32-1:0] _mystream_a2_source_fsm_2;
  localparam _mystream_a2_source_fsm_2_init = 0;
  wire _set_flag_194;
  assign _set_flag_194 = th_comp == 17;
  assign ram_a_3_0_addr = (_mystream_stream_oready && _mystream_a3_source_ram_renable && (_mystream_a3_source_sel == 4))? _mystream_a3_source_ram_raddr : 
                          ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_addr_49 : 'hx;
  assign ram_a_3_0_enable = (_mystream_stream_oready && _mystream_a3_source_ram_renable && (_mystream_a3_source_sel == 4))? 1'd1 : 
                            ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  localparam _tmp_195 = 1;
  wire [_tmp_195-1:0] _tmp_196;
  assign _tmp_196 = _mystream_stream_oready && _mystream_a3_source_ram_renable && (_mystream_a3_source_sel == 4);
  reg [_tmp_195-1:0] __tmp_196_1;
  assign _mystream_a3_source_ram_rdata = (_mystream_a3_source_sel == 4)? ram_a_3_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_5;
  assign mystream_a3_data = __variable_wdata_5;
  reg [32-1:0] _mystream_a3_source_fsm_3;
  localparam _mystream_a3_source_fsm_3_init = 0;
  wire _set_flag_197;
  assign _set_flag_197 = th_comp == 18;
  assign ram_a_4_0_addr = (_mystream_stream_oready && _mystream_a4_source_ram_renable && (_mystream_a4_source_sel == 5))? _mystream_a4_source_ram_raddr : 
                          ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_addr_51 : 'hx;
  assign ram_a_4_0_enable = (_mystream_stream_oready && _mystream_a4_source_ram_renable && (_mystream_a4_source_sel == 5))? 1'd1 : 
                            ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  localparam _tmp_198 = 1;
  wire [_tmp_198-1:0] _tmp_199;
  assign _tmp_199 = _mystream_stream_oready && _mystream_a4_source_ram_renable && (_mystream_a4_source_sel == 5);
  reg [_tmp_198-1:0] __tmp_199_1;
  assign _mystream_a4_source_ram_rdata = (_mystream_a4_source_sel == 5)? ram_a_4_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_6;
  assign mystream_a4_data = __variable_wdata_6;
  reg [32-1:0] _mystream_a4_source_fsm_4;
  localparam _mystream_a4_source_fsm_4_init = 0;
  wire _set_flag_200;
  assign _set_flag_200 = th_comp == 19;
  assign ram_a_5_0_addr = (_mystream_stream_oready && _mystream_a5_source_ram_renable && (_mystream_a5_source_sel == 6))? _mystream_a5_source_ram_raddr : 
                          ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_addr_53 : 'hx;
  assign ram_a_5_0_enable = (_mystream_stream_oready && _mystream_a5_source_ram_renable && (_mystream_a5_source_sel == 6))? 1'd1 : 
                            ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  localparam _tmp_201 = 1;
  wire [_tmp_201-1:0] _tmp_202;
  assign _tmp_202 = _mystream_stream_oready && _mystream_a5_source_ram_renable && (_mystream_a5_source_sel == 6);
  reg [_tmp_201-1:0] __tmp_202_1;
  assign _mystream_a5_source_ram_rdata = (_mystream_a5_source_sel == 6)? ram_a_5_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_7;
  assign mystream_a5_data = __variable_wdata_7;
  reg [32-1:0] _mystream_a5_source_fsm_5;
  localparam _mystream_a5_source_fsm_5_init = 0;
  wire _set_flag_203;
  assign _set_flag_203 = th_comp == 20;
  assign ram_a_6_0_addr = (_mystream_stream_oready && _mystream_a6_source_ram_renable && (_mystream_a6_source_sel == 7))? _mystream_a6_source_ram_raddr : 
                          ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_addr_55 : 'hx;
  assign ram_a_6_0_enable = (_mystream_stream_oready && _mystream_a6_source_ram_renable && (_mystream_a6_source_sel == 7))? 1'd1 : 
                            ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  localparam _tmp_204 = 1;
  wire [_tmp_204-1:0] _tmp_205;
  assign _tmp_205 = _mystream_stream_oready && _mystream_a6_source_ram_renable && (_mystream_a6_source_sel == 7);
  reg [_tmp_204-1:0] __tmp_205_1;
  assign _mystream_a6_source_ram_rdata = (_mystream_a6_source_sel == 7)? ram_a_6_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_8;
  assign mystream_a6_data = __variable_wdata_8;
  reg [32-1:0] _mystream_a6_source_fsm_6;
  localparam _mystream_a6_source_fsm_6_init = 0;
  wire _set_flag_206;
  assign _set_flag_206 = th_comp == 21;
  assign ram_a_7_0_addr = (_mystream_stream_oready && _mystream_a7_source_ram_renable && (_mystream_a7_source_sel == 8))? _mystream_a7_source_ram_raddr : 
                          ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_addr_57 : 'hx;
  assign ram_a_7_0_enable = (_mystream_stream_oready && _mystream_a7_source_ram_renable && (_mystream_a7_source_sel == 8))? 1'd1 : 
                            ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  localparam _tmp_207 = 1;
  wire [_tmp_207-1:0] _tmp_208;
  assign _tmp_208 = _mystream_stream_oready && _mystream_a7_source_ram_renable && (_mystream_a7_source_sel == 8);
  reg [_tmp_207-1:0] __tmp_208_1;
  assign _mystream_a7_source_ram_rdata = (_mystream_a7_source_sel == 8)? ram_a_7_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_9;
  assign mystream_a7_data = __variable_wdata_9;
  reg [32-1:0] _mystream_a7_source_fsm_7;
  localparam _mystream_a7_source_fsm_7_init = 0;
  wire _set_flag_209;
  assign _set_flag_209 = th_comp == 22;
  assign ram_a_8_0_addr = (_mystream_stream_oready && _mystream_a8_source_ram_renable && (_mystream_a8_source_sel == 9))? _mystream_a8_source_ram_raddr : 
                          ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_addr_59 : 'hx;
  assign ram_a_8_0_enable = (_mystream_stream_oready && _mystream_a8_source_ram_renable && (_mystream_a8_source_sel == 9))? 1'd1 : 
                            ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  localparam _tmp_210 = 1;
  wire [_tmp_210-1:0] _tmp_211;
  assign _tmp_211 = _mystream_stream_oready && _mystream_a8_source_ram_renable && (_mystream_a8_source_sel == 9);
  reg [_tmp_210-1:0] __tmp_211_1;
  assign _mystream_a8_source_ram_rdata = (_mystream_a8_source_sel == 9)? ram_a_8_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_10;
  assign mystream_a8_data = __variable_wdata_10;
  reg [32-1:0] _mystream_a8_source_fsm_8;
  localparam _mystream_a8_source_fsm_8_init = 0;
  wire _set_flag_212;
  assign _set_flag_212 = th_comp == 23;
  assign ram_a_9_0_addr = (_mystream_stream_oready && _mystream_a9_source_ram_renable && (_mystream_a9_source_sel == 10))? _mystream_a9_source_ram_raddr : 
                          ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_addr_61 : 'hx;
  assign ram_a_9_0_enable = (_mystream_stream_oready && _mystream_a9_source_ram_renable && (_mystream_a9_source_sel == 10))? 1'd1 : 
                            ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  localparam _tmp_213 = 1;
  wire [_tmp_213-1:0] _tmp_214;
  assign _tmp_214 = _mystream_stream_oready && _mystream_a9_source_ram_renable && (_mystream_a9_source_sel == 10);
  reg [_tmp_213-1:0] __tmp_214_1;
  assign _mystream_a9_source_ram_rdata = (_mystream_a9_source_sel == 10)? ram_a_9_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_11;
  assign mystream_a9_data = __variable_wdata_11;
  reg [32-1:0] _mystream_a9_source_fsm_9;
  localparam _mystream_a9_source_fsm_9_init = 0;
  wire _set_flag_215;
  assign _set_flag_215 = th_comp == 24;
  assign ram_a_10_0_addr = (_mystream_stream_oready && _mystream_a10_source_ram_renable && (_mystream_a10_source_sel == 11))? _mystream_a10_source_ram_raddr : 
                           ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_addr_63 : 'hx;
  assign ram_a_10_0_enable = (_mystream_stream_oready && _mystream_a10_source_ram_renable && (_mystream_a10_source_sel == 11))? 1'd1 : 
                             ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  localparam _tmp_216 = 1;
  wire [_tmp_216-1:0] _tmp_217;
  assign _tmp_217 = _mystream_stream_oready && _mystream_a10_source_ram_renable && (_mystream_a10_source_sel == 11);
  reg [_tmp_216-1:0] __tmp_217_1;
  assign _mystream_a10_source_ram_rdata = (_mystream_a10_source_sel == 11)? ram_a_10_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_12;
  assign mystream_a10_data = __variable_wdata_12;
  reg [32-1:0] _mystream_a10_source_fsm_10;
  localparam _mystream_a10_source_fsm_10_init = 0;
  wire _set_flag_218;
  assign _set_flag_218 = th_comp == 25;
  assign ram_a_11_0_addr = (_mystream_stream_oready && _mystream_a11_source_ram_renable && (_mystream_a11_source_sel == 12))? _mystream_a11_source_ram_raddr : 
                           ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_addr_65 : 'hx;
  assign ram_a_11_0_enable = (_mystream_stream_oready && _mystream_a11_source_ram_renable && (_mystream_a11_source_sel == 12))? 1'd1 : 
                             ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  localparam _tmp_219 = 1;
  wire [_tmp_219-1:0] _tmp_220;
  assign _tmp_220 = _mystream_stream_oready && _mystream_a11_source_ram_renable && (_mystream_a11_source_sel == 12);
  reg [_tmp_219-1:0] __tmp_220_1;
  assign _mystream_a11_source_ram_rdata = (_mystream_a11_source_sel == 12)? ram_a_11_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_13;
  assign mystream_a11_data = __variable_wdata_13;
  reg [32-1:0] _mystream_a11_source_fsm_11;
  localparam _mystream_a11_source_fsm_11_init = 0;
  wire _set_flag_221;
  assign _set_flag_221 = th_comp == 26;
  assign ram_a_12_0_addr = (_mystream_stream_oready && _mystream_a12_source_ram_renable && (_mystream_a12_source_sel == 13))? _mystream_a12_source_ram_raddr : 
                           ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_addr_67 : 'hx;
  assign ram_a_12_0_enable = (_mystream_stream_oready && _mystream_a12_source_ram_renable && (_mystream_a12_source_sel == 13))? 1'd1 : 
                             ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  localparam _tmp_222 = 1;
  wire [_tmp_222-1:0] _tmp_223;
  assign _tmp_223 = _mystream_stream_oready && _mystream_a12_source_ram_renable && (_mystream_a12_source_sel == 13);
  reg [_tmp_222-1:0] __tmp_223_1;
  assign _mystream_a12_source_ram_rdata = (_mystream_a12_source_sel == 13)? ram_a_12_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_14;
  assign mystream_a12_data = __variable_wdata_14;
  reg [32-1:0] _mystream_a12_source_fsm_12;
  localparam _mystream_a12_source_fsm_12_init = 0;
  wire _set_flag_224;
  assign _set_flag_224 = th_comp == 27;
  assign ram_a_13_0_addr = (_mystream_stream_oready && _mystream_a13_source_ram_renable && (_mystream_a13_source_sel == 14))? _mystream_a13_source_ram_raddr : 
                           ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_addr_69 : 'hx;
  assign ram_a_13_0_enable = (_mystream_stream_oready && _mystream_a13_source_ram_renable && (_mystream_a13_source_sel == 14))? 1'd1 : 
                             ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  localparam _tmp_225 = 1;
  wire [_tmp_225-1:0] _tmp_226;
  assign _tmp_226 = _mystream_stream_oready && _mystream_a13_source_ram_renable && (_mystream_a13_source_sel == 14);
  reg [_tmp_225-1:0] __tmp_226_1;
  assign _mystream_a13_source_ram_rdata = (_mystream_a13_source_sel == 14)? ram_a_13_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_15;
  assign mystream_a13_data = __variable_wdata_15;
  reg [32-1:0] _mystream_a13_source_fsm_13;
  localparam _mystream_a13_source_fsm_13_init = 0;
  wire _set_flag_227;
  assign _set_flag_227 = th_comp == 28;
  assign ram_a_14_0_addr = (_mystream_stream_oready && _mystream_a14_source_ram_renable && (_mystream_a14_source_sel == 15))? _mystream_a14_source_ram_raddr : 
                           ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_addr_71 : 'hx;
  assign ram_a_14_0_enable = (_mystream_stream_oready && _mystream_a14_source_ram_renable && (_mystream_a14_source_sel == 15))? 1'd1 : 
                             ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  localparam _tmp_228 = 1;
  wire [_tmp_228-1:0] _tmp_229;
  assign _tmp_229 = _mystream_stream_oready && _mystream_a14_source_ram_renable && (_mystream_a14_source_sel == 15);
  reg [_tmp_228-1:0] __tmp_229_1;
  assign _mystream_a14_source_ram_rdata = (_mystream_a14_source_sel == 15)? ram_a_14_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_16;
  assign mystream_a14_data = __variable_wdata_16;
  reg [32-1:0] _mystream_a14_source_fsm_14;
  localparam _mystream_a14_source_fsm_14_init = 0;
  wire _set_flag_230;
  assign _set_flag_230 = th_comp == 29;
  assign ram_a_15_0_addr = (_mystream_stream_oready && _mystream_a15_source_ram_renable && (_mystream_a15_source_sel == 16))? _mystream_a15_source_ram_raddr : 
                           ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_addr_73 : 'hx;
  assign ram_a_15_0_enable = (_mystream_stream_oready && _mystream_a15_source_ram_renable && (_mystream_a15_source_sel == 16))? 1'd1 : 
                             ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  localparam _tmp_231 = 1;
  wire [_tmp_231-1:0] _tmp_232;
  assign _tmp_232 = _mystream_stream_oready && _mystream_a15_source_ram_renable && (_mystream_a15_source_sel == 16);
  reg [_tmp_231-1:0] __tmp_232_1;
  assign _mystream_a15_source_ram_rdata = (_mystream_a15_source_sel == 16)? ram_a_15_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_17;
  assign mystream_a15_data = __variable_wdata_17;
  reg [32-1:0] _mystream_a15_source_fsm_15;
  localparam _mystream_a15_source_fsm_15_init = 0;
  wire _set_flag_233;
  assign _set_flag_233 = th_comp == 30;
  assign ram_a_16_0_addr = (_mystream_stream_oready && _mystream_a16_source_ram_renable && (_mystream_a16_source_sel == 17))? _mystream_a16_source_ram_raddr : 
                           ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_addr_75 : 'hx;
  assign ram_a_16_0_enable = (_mystream_stream_oready && _mystream_a16_source_ram_renable && (_mystream_a16_source_sel == 17))? 1'd1 : 
                             ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  localparam _tmp_234 = 1;
  wire [_tmp_234-1:0] _tmp_235;
  assign _tmp_235 = _mystream_stream_oready && _mystream_a16_source_ram_renable && (_mystream_a16_source_sel == 17);
  reg [_tmp_234-1:0] __tmp_235_1;
  assign _mystream_a16_source_ram_rdata = (_mystream_a16_source_sel == 17)? ram_a_16_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_18;
  assign mystream_a16_data = __variable_wdata_18;
  reg [32-1:0] _mystream_a16_source_fsm_16;
  localparam _mystream_a16_source_fsm_16_init = 0;
  wire _set_flag_236;
  assign _set_flag_236 = th_comp == 31;
  assign ram_a_17_0_addr = (_mystream_stream_oready && _mystream_a17_source_ram_renable && (_mystream_a17_source_sel == 18))? _mystream_a17_source_ram_raddr : 
                           ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_addr_77 : 'hx;
  assign ram_a_17_0_enable = (_mystream_stream_oready && _mystream_a17_source_ram_renable && (_mystream_a17_source_sel == 18))? 1'd1 : 
                             ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  localparam _tmp_237 = 1;
  wire [_tmp_237-1:0] _tmp_238;
  assign _tmp_238 = _mystream_stream_oready && _mystream_a17_source_ram_renable && (_mystream_a17_source_sel == 18);
  reg [_tmp_237-1:0] __tmp_238_1;
  assign _mystream_a17_source_ram_rdata = (_mystream_a17_source_sel == 18)? ram_a_17_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_19;
  assign mystream_a17_data = __variable_wdata_19;
  reg [32-1:0] _mystream_a17_source_fsm_17;
  localparam _mystream_a17_source_fsm_17_init = 0;
  wire _set_flag_239;
  assign _set_flag_239 = th_comp == 32;
  assign ram_a_18_0_addr = (_mystream_stream_oready && _mystream_a18_source_ram_renable && (_mystream_a18_source_sel == 19))? _mystream_a18_source_ram_raddr : 
                           ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_addr_79 : 'hx;
  assign ram_a_18_0_enable = (_mystream_stream_oready && _mystream_a18_source_ram_renable && (_mystream_a18_source_sel == 19))? 1'd1 : 
                             ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  localparam _tmp_240 = 1;
  wire [_tmp_240-1:0] _tmp_241;
  assign _tmp_241 = _mystream_stream_oready && _mystream_a18_source_ram_renable && (_mystream_a18_source_sel == 19);
  reg [_tmp_240-1:0] __tmp_241_1;
  assign _mystream_a18_source_ram_rdata = (_mystream_a18_source_sel == 19)? ram_a_18_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_20;
  assign mystream_a18_data = __variable_wdata_20;
  reg [32-1:0] _mystream_a18_source_fsm_18;
  localparam _mystream_a18_source_fsm_18_init = 0;
  wire _set_flag_242;
  assign _set_flag_242 = th_comp == 33;
  assign ram_a_19_0_addr = (_mystream_stream_oready && _mystream_a19_source_ram_renable && (_mystream_a19_source_sel == 20))? _mystream_a19_source_ram_raddr : 
                           ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_addr_81 : 'hx;
  assign ram_a_19_0_enable = (_mystream_stream_oready && _mystream_a19_source_ram_renable && (_mystream_a19_source_sel == 20))? 1'd1 : 
                             ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  localparam _tmp_243 = 1;
  wire [_tmp_243-1:0] _tmp_244;
  assign _tmp_244 = _mystream_stream_oready && _mystream_a19_source_ram_renable && (_mystream_a19_source_sel == 20);
  reg [_tmp_243-1:0] __tmp_244_1;
  assign _mystream_a19_source_ram_rdata = (_mystream_a19_source_sel == 20)? ram_a_19_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_21;
  assign mystream_a19_data = __variable_wdata_21;
  reg [32-1:0] _mystream_a19_source_fsm_19;
  localparam _mystream_a19_source_fsm_19_init = 0;
  wire _set_flag_245;
  assign _set_flag_245 = th_comp == 34;
  assign ram_a_20_0_addr = (_mystream_stream_oready && _mystream_a20_source_ram_renable && (_mystream_a20_source_sel == 21))? _mystream_a20_source_ram_raddr : 
                           ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_addr_83 : 'hx;
  assign ram_a_20_0_enable = (_mystream_stream_oready && _mystream_a20_source_ram_renable && (_mystream_a20_source_sel == 21))? 1'd1 : 
                             ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  localparam _tmp_246 = 1;
  wire [_tmp_246-1:0] _tmp_247;
  assign _tmp_247 = _mystream_stream_oready && _mystream_a20_source_ram_renable && (_mystream_a20_source_sel == 21);
  reg [_tmp_246-1:0] __tmp_247_1;
  assign _mystream_a20_source_ram_rdata = (_mystream_a20_source_sel == 21)? ram_a_20_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_22;
  assign mystream_a20_data = __variable_wdata_22;
  reg [32-1:0] _mystream_a20_source_fsm_20;
  localparam _mystream_a20_source_fsm_20_init = 0;
  wire _set_flag_248;
  assign _set_flag_248 = th_comp == 35;
  assign ram_a_21_0_addr = (_mystream_stream_oready && _mystream_a21_source_ram_renable && (_mystream_a21_source_sel == 22))? _mystream_a21_source_ram_raddr : 
                           ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_addr_85 : 'hx;
  assign ram_a_21_0_enable = (_mystream_stream_oready && _mystream_a21_source_ram_renable && (_mystream_a21_source_sel == 22))? 1'd1 : 
                             ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  localparam _tmp_249 = 1;
  wire [_tmp_249-1:0] _tmp_250;
  assign _tmp_250 = _mystream_stream_oready && _mystream_a21_source_ram_renable && (_mystream_a21_source_sel == 22);
  reg [_tmp_249-1:0] __tmp_250_1;
  assign _mystream_a21_source_ram_rdata = (_mystream_a21_source_sel == 22)? ram_a_21_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_23;
  assign mystream_a21_data = __variable_wdata_23;
  reg [32-1:0] _mystream_a21_source_fsm_21;
  localparam _mystream_a21_source_fsm_21_init = 0;
  wire _set_flag_251;
  assign _set_flag_251 = th_comp == 36;
  assign ram_a_22_0_addr = (_mystream_stream_oready && _mystream_a22_source_ram_renable && (_mystream_a22_source_sel == 23))? _mystream_a22_source_ram_raddr : 
                           ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_addr_87 : 'hx;
  assign ram_a_22_0_enable = (_mystream_stream_oready && _mystream_a22_source_ram_renable && (_mystream_a22_source_sel == 23))? 1'd1 : 
                             ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  localparam _tmp_252 = 1;
  wire [_tmp_252-1:0] _tmp_253;
  assign _tmp_253 = _mystream_stream_oready && _mystream_a22_source_ram_renable && (_mystream_a22_source_sel == 23);
  reg [_tmp_252-1:0] __tmp_253_1;
  assign _mystream_a22_source_ram_rdata = (_mystream_a22_source_sel == 23)? ram_a_22_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_24;
  assign mystream_a22_data = __variable_wdata_24;
  reg [32-1:0] _mystream_a22_source_fsm_22;
  localparam _mystream_a22_source_fsm_22_init = 0;
  wire _set_flag_254;
  assign _set_flag_254 = th_comp == 37;
  assign ram_a_23_0_addr = (_mystream_stream_oready && _mystream_a23_source_ram_renable && (_mystream_a23_source_sel == 24))? _mystream_a23_source_ram_raddr : 
                           ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_addr_89 : 'hx;
  assign ram_a_23_0_enable = (_mystream_stream_oready && _mystream_a23_source_ram_renable && (_mystream_a23_source_sel == 24))? 1'd1 : 
                             ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  localparam _tmp_255 = 1;
  wire [_tmp_255-1:0] _tmp_256;
  assign _tmp_256 = _mystream_stream_oready && _mystream_a23_source_ram_renable && (_mystream_a23_source_sel == 24);
  reg [_tmp_255-1:0] __tmp_256_1;
  assign _mystream_a23_source_ram_rdata = (_mystream_a23_source_sel == 24)? ram_a_23_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_25;
  assign mystream_a23_data = __variable_wdata_25;
  reg [32-1:0] _mystream_a23_source_fsm_23;
  localparam _mystream_a23_source_fsm_23_init = 0;
  wire _set_flag_257;
  assign _set_flag_257 = th_comp == 38;
  assign ram_a_24_0_addr = (_mystream_stream_oready && _mystream_a24_source_ram_renable && (_mystream_a24_source_sel == 25))? _mystream_a24_source_ram_raddr : 
                           ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_addr_91 : 'hx;
  assign ram_a_24_0_enable = (_mystream_stream_oready && _mystream_a24_source_ram_renable && (_mystream_a24_source_sel == 25))? 1'd1 : 
                             ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  localparam _tmp_258 = 1;
  wire [_tmp_258-1:0] _tmp_259;
  assign _tmp_259 = _mystream_stream_oready && _mystream_a24_source_ram_renable && (_mystream_a24_source_sel == 25);
  reg [_tmp_258-1:0] __tmp_259_1;
  assign _mystream_a24_source_ram_rdata = (_mystream_a24_source_sel == 25)? ram_a_24_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_26;
  assign mystream_a24_data = __variable_wdata_26;
  reg [32-1:0] _mystream_a24_source_fsm_24;
  localparam _mystream_a24_source_fsm_24_init = 0;
  wire _set_flag_260;
  assign _set_flag_260 = th_comp == 39;
  assign ram_a_25_0_addr = (_mystream_stream_oready && _mystream_a25_source_ram_renable && (_mystream_a25_source_sel == 26))? _mystream_a25_source_ram_raddr : 
                           ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_addr_93 : 'hx;
  assign ram_a_25_0_enable = (_mystream_stream_oready && _mystream_a25_source_ram_renable && (_mystream_a25_source_sel == 26))? 1'd1 : 
                             ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  localparam _tmp_261 = 1;
  wire [_tmp_261-1:0] _tmp_262;
  assign _tmp_262 = _mystream_stream_oready && _mystream_a25_source_ram_renable && (_mystream_a25_source_sel == 26);
  reg [_tmp_261-1:0] __tmp_262_1;
  assign _mystream_a25_source_ram_rdata = (_mystream_a25_source_sel == 26)? ram_a_25_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_27;
  assign mystream_a25_data = __variable_wdata_27;
  reg [32-1:0] _mystream_a25_source_fsm_25;
  localparam _mystream_a25_source_fsm_25_init = 0;
  wire _set_flag_263;
  assign _set_flag_263 = th_comp == 40;
  assign ram_a_26_0_addr = (_mystream_stream_oready && _mystream_a26_source_ram_renable && (_mystream_a26_source_sel == 27))? _mystream_a26_source_ram_raddr : 
                           ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_addr_95 : 'hx;
  assign ram_a_26_0_enable = (_mystream_stream_oready && _mystream_a26_source_ram_renable && (_mystream_a26_source_sel == 27))? 1'd1 : 
                             ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  localparam _tmp_264 = 1;
  wire [_tmp_264-1:0] _tmp_265;
  assign _tmp_265 = _mystream_stream_oready && _mystream_a26_source_ram_renable && (_mystream_a26_source_sel == 27);
  reg [_tmp_264-1:0] __tmp_265_1;
  assign _mystream_a26_source_ram_rdata = (_mystream_a26_source_sel == 27)? ram_a_26_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_28;
  assign mystream_a26_data = __variable_wdata_28;
  reg [32-1:0] _mystream_a26_source_fsm_26;
  localparam _mystream_a26_source_fsm_26_init = 0;
  wire _set_flag_266;
  assign _set_flag_266 = th_comp == 41;
  assign ram_a_27_0_addr = (_mystream_stream_oready && _mystream_a27_source_ram_renable && (_mystream_a27_source_sel == 28))? _mystream_a27_source_ram_raddr : 
                           ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_addr_97 : 'hx;
  assign ram_a_27_0_enable = (_mystream_stream_oready && _mystream_a27_source_ram_renable && (_mystream_a27_source_sel == 28))? 1'd1 : 
                             ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  localparam _tmp_267 = 1;
  wire [_tmp_267-1:0] _tmp_268;
  assign _tmp_268 = _mystream_stream_oready && _mystream_a27_source_ram_renable && (_mystream_a27_source_sel == 28);
  reg [_tmp_267-1:0] __tmp_268_1;
  assign _mystream_a27_source_ram_rdata = (_mystream_a27_source_sel == 28)? ram_a_27_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_29;
  assign mystream_a27_data = __variable_wdata_29;
  reg [32-1:0] _mystream_a27_source_fsm_27;
  localparam _mystream_a27_source_fsm_27_init = 0;
  wire _set_flag_269;
  assign _set_flag_269 = th_comp == 42;
  assign ram_a_28_0_addr = (_mystream_stream_oready && _mystream_a28_source_ram_renable && (_mystream_a28_source_sel == 29))? _mystream_a28_source_ram_raddr : 
                           ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_addr_99 : 'hx;
  assign ram_a_28_0_enable = (_mystream_stream_oready && _mystream_a28_source_ram_renable && (_mystream_a28_source_sel == 29))? 1'd1 : 
                             ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  localparam _tmp_270 = 1;
  wire [_tmp_270-1:0] _tmp_271;
  assign _tmp_271 = _mystream_stream_oready && _mystream_a28_source_ram_renable && (_mystream_a28_source_sel == 29);
  reg [_tmp_270-1:0] __tmp_271_1;
  assign _mystream_a28_source_ram_rdata = (_mystream_a28_source_sel == 29)? ram_a_28_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_30;
  assign mystream_a28_data = __variable_wdata_30;
  reg [32-1:0] _mystream_a28_source_fsm_28;
  localparam _mystream_a28_source_fsm_28_init = 0;
  wire _set_flag_272;
  assign _set_flag_272 = th_comp == 43;
  assign ram_a_29_0_addr = (_mystream_stream_oready && _mystream_a29_source_ram_renable && (_mystream_a29_source_sel == 30))? _mystream_a29_source_ram_raddr : 
                           ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_addr_101 : 'hx;
  assign ram_a_29_0_enable = (_mystream_stream_oready && _mystream_a29_source_ram_renable && (_mystream_a29_source_sel == 30))? 1'd1 : 
                             ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  localparam _tmp_273 = 1;
  wire [_tmp_273-1:0] _tmp_274;
  assign _tmp_274 = _mystream_stream_oready && _mystream_a29_source_ram_renable && (_mystream_a29_source_sel == 30);
  reg [_tmp_273-1:0] __tmp_274_1;
  assign _mystream_a29_source_ram_rdata = (_mystream_a29_source_sel == 30)? ram_a_29_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_31;
  assign mystream_a29_data = __variable_wdata_31;
  reg [32-1:0] _mystream_a29_source_fsm_29;
  localparam _mystream_a29_source_fsm_29_init = 0;
  wire _set_flag_275;
  assign _set_flag_275 = th_comp == 44;
  assign ram_a_30_0_addr = (_mystream_stream_oready && _mystream_a30_source_ram_renable && (_mystream_a30_source_sel == 31))? _mystream_a30_source_ram_raddr : 
                           ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_addr_103 : 'hx;
  assign ram_a_30_0_enable = (_mystream_stream_oready && _mystream_a30_source_ram_renable && (_mystream_a30_source_sel == 31))? 1'd1 : 
                             ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  localparam _tmp_276 = 1;
  wire [_tmp_276-1:0] _tmp_277;
  assign _tmp_277 = _mystream_stream_oready && _mystream_a30_source_ram_renable && (_mystream_a30_source_sel == 31);
  reg [_tmp_276-1:0] __tmp_277_1;
  assign _mystream_a30_source_ram_rdata = (_mystream_a30_source_sel == 31)? ram_a_30_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_32;
  assign mystream_a30_data = __variable_wdata_32;
  reg [32-1:0] _mystream_a30_source_fsm_30;
  localparam _mystream_a30_source_fsm_30_init = 0;
  wire _set_flag_278;
  assign _set_flag_278 = th_comp == 45;
  assign ram_a_31_0_addr = (_mystream_stream_oready && _mystream_a31_source_ram_renable && (_mystream_a31_source_sel == 32))? _mystream_a31_source_ram_raddr : 
                           ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? write_burst_packed_ram_addr_105 : 'hx;
  assign ram_a_31_0_enable = (_mystream_stream_oready && _mystream_a31_source_ram_renable && (_mystream_a31_source_sel == 32))? 1'd1 : 
                             ((write_burst_packed_fsm_0 == 1) && _myaxi_read_narrow_wvalid_37)? 1'd1 : 0;
  localparam _tmp_279 = 1;
  wire [_tmp_279-1:0] _tmp_280;
  assign _tmp_280 = _mystream_stream_oready && _mystream_a31_source_ram_renable && (_mystream_a31_source_sel == 32);
  reg [_tmp_279-1:0] __tmp_280_1;
  assign _mystream_a31_source_ram_rdata = (_mystream_a31_source_sel == 32)? ram_a_31_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_33;
  assign mystream_a31_data = __variable_wdata_33;
  reg [32-1:0] _mystream_a31_source_fsm_31;
  localparam _mystream_a31_source_fsm_31_init = 0;
  wire _set_flag_281;
  assign _set_flag_281 = th_comp == 48;
  assign ram_b_0_0_addr = (_mystream_stream_oready && _mystream_b0_source_ram_renable && (_mystream_b0_source_sel == 33))? _mystream_b0_source_ram_raddr : 
                          ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_addr_119 : 'hx;
  assign ram_b_0_0_enable = (_mystream_stream_oready && _mystream_b0_source_ram_renable && (_mystream_b0_source_sel == 33))? 1'd1 : 
                            ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  localparam _tmp_282 = 1;
  wire [_tmp_282-1:0] _tmp_283;
  assign _tmp_283 = _mystream_stream_oready && _mystream_b0_source_ram_renable && (_mystream_b0_source_sel == 33);
  reg [_tmp_282-1:0] __tmp_283_1;
  assign _mystream_b0_source_ram_rdata = (_mystream_b0_source_sel == 33)? ram_b_0_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_34;
  assign mystream_b0_data = __variable_wdata_34;
  reg [32-1:0] _mystream_b0_source_fsm_32;
  localparam _mystream_b0_source_fsm_32_init = 0;
  wire _set_flag_284;
  assign _set_flag_284 = th_comp == 49;
  assign ram_b_1_0_addr = (_mystream_stream_oready && _mystream_b1_source_ram_renable && (_mystream_b1_source_sel == 34))? _mystream_b1_source_ram_raddr : 
                          ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_addr_121 : 'hx;
  assign ram_b_1_0_enable = (_mystream_stream_oready && _mystream_b1_source_ram_renable && (_mystream_b1_source_sel == 34))? 1'd1 : 
                            ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  localparam _tmp_285 = 1;
  wire [_tmp_285-1:0] _tmp_286;
  assign _tmp_286 = _mystream_stream_oready && _mystream_b1_source_ram_renable && (_mystream_b1_source_sel == 34);
  reg [_tmp_285-1:0] __tmp_286_1;
  assign _mystream_b1_source_ram_rdata = (_mystream_b1_source_sel == 34)? ram_b_1_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_35;
  assign mystream_b1_data = __variable_wdata_35;
  reg [32-1:0] _mystream_b1_source_fsm_33;
  localparam _mystream_b1_source_fsm_33_init = 0;
  wire _set_flag_287;
  assign _set_flag_287 = th_comp == 50;
  assign ram_b_2_0_addr = (_mystream_stream_oready && _mystream_b2_source_ram_renable && (_mystream_b2_source_sel == 35))? _mystream_b2_source_ram_raddr : 
                          ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_addr_123 : 'hx;
  assign ram_b_2_0_enable = (_mystream_stream_oready && _mystream_b2_source_ram_renable && (_mystream_b2_source_sel == 35))? 1'd1 : 
                            ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  localparam _tmp_288 = 1;
  wire [_tmp_288-1:0] _tmp_289;
  assign _tmp_289 = _mystream_stream_oready && _mystream_b2_source_ram_renable && (_mystream_b2_source_sel == 35);
  reg [_tmp_288-1:0] __tmp_289_1;
  assign _mystream_b2_source_ram_rdata = (_mystream_b2_source_sel == 35)? ram_b_2_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_36;
  assign mystream_b2_data = __variable_wdata_36;
  reg [32-1:0] _mystream_b2_source_fsm_34;
  localparam _mystream_b2_source_fsm_34_init = 0;
  wire _set_flag_290;
  assign _set_flag_290 = th_comp == 51;
  assign ram_b_3_0_addr = (_mystream_stream_oready && _mystream_b3_source_ram_renable && (_mystream_b3_source_sel == 36))? _mystream_b3_source_ram_raddr : 
                          ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_addr_125 : 'hx;
  assign ram_b_3_0_enable = (_mystream_stream_oready && _mystream_b3_source_ram_renable && (_mystream_b3_source_sel == 36))? 1'd1 : 
                            ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  localparam _tmp_291 = 1;
  wire [_tmp_291-1:0] _tmp_292;
  assign _tmp_292 = _mystream_stream_oready && _mystream_b3_source_ram_renable && (_mystream_b3_source_sel == 36);
  reg [_tmp_291-1:0] __tmp_292_1;
  assign _mystream_b3_source_ram_rdata = (_mystream_b3_source_sel == 36)? ram_b_3_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_37;
  assign mystream_b3_data = __variable_wdata_37;
  reg [32-1:0] _mystream_b3_source_fsm_35;
  localparam _mystream_b3_source_fsm_35_init = 0;
  wire _set_flag_293;
  assign _set_flag_293 = th_comp == 52;
  assign ram_b_4_0_addr = (_mystream_stream_oready && _mystream_b4_source_ram_renable && (_mystream_b4_source_sel == 37))? _mystream_b4_source_ram_raddr : 
                          ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_addr_127 : 'hx;
  assign ram_b_4_0_enable = (_mystream_stream_oready && _mystream_b4_source_ram_renable && (_mystream_b4_source_sel == 37))? 1'd1 : 
                            ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  localparam _tmp_294 = 1;
  wire [_tmp_294-1:0] _tmp_295;
  assign _tmp_295 = _mystream_stream_oready && _mystream_b4_source_ram_renable && (_mystream_b4_source_sel == 37);
  reg [_tmp_294-1:0] __tmp_295_1;
  assign _mystream_b4_source_ram_rdata = (_mystream_b4_source_sel == 37)? ram_b_4_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_38;
  assign mystream_b4_data = __variable_wdata_38;
  reg [32-1:0] _mystream_b4_source_fsm_36;
  localparam _mystream_b4_source_fsm_36_init = 0;
  wire _set_flag_296;
  assign _set_flag_296 = th_comp == 53;
  assign ram_b_5_0_addr = (_mystream_stream_oready && _mystream_b5_source_ram_renable && (_mystream_b5_source_sel == 38))? _mystream_b5_source_ram_raddr : 
                          ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_addr_129 : 'hx;
  assign ram_b_5_0_enable = (_mystream_stream_oready && _mystream_b5_source_ram_renable && (_mystream_b5_source_sel == 38))? 1'd1 : 
                            ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  localparam _tmp_297 = 1;
  wire [_tmp_297-1:0] _tmp_298;
  assign _tmp_298 = _mystream_stream_oready && _mystream_b5_source_ram_renable && (_mystream_b5_source_sel == 38);
  reg [_tmp_297-1:0] __tmp_298_1;
  assign _mystream_b5_source_ram_rdata = (_mystream_b5_source_sel == 38)? ram_b_5_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_39;
  assign mystream_b5_data = __variable_wdata_39;
  reg [32-1:0] _mystream_b5_source_fsm_37;
  localparam _mystream_b5_source_fsm_37_init = 0;
  wire _set_flag_299;
  assign _set_flag_299 = th_comp == 54;
  assign ram_b_6_0_addr = (_mystream_stream_oready && _mystream_b6_source_ram_renable && (_mystream_b6_source_sel == 39))? _mystream_b6_source_ram_raddr : 
                          ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_addr_131 : 'hx;
  assign ram_b_6_0_enable = (_mystream_stream_oready && _mystream_b6_source_ram_renable && (_mystream_b6_source_sel == 39))? 1'd1 : 
                            ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  localparam _tmp_300 = 1;
  wire [_tmp_300-1:0] _tmp_301;
  assign _tmp_301 = _mystream_stream_oready && _mystream_b6_source_ram_renable && (_mystream_b6_source_sel == 39);
  reg [_tmp_300-1:0] __tmp_301_1;
  assign _mystream_b6_source_ram_rdata = (_mystream_b6_source_sel == 39)? ram_b_6_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_40;
  assign mystream_b6_data = __variable_wdata_40;
  reg [32-1:0] _mystream_b6_source_fsm_38;
  localparam _mystream_b6_source_fsm_38_init = 0;
  wire _set_flag_302;
  assign _set_flag_302 = th_comp == 55;
  assign ram_b_7_0_addr = (_mystream_stream_oready && _mystream_b7_source_ram_renable && (_mystream_b7_source_sel == 40))? _mystream_b7_source_ram_raddr : 
                          ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_addr_133 : 'hx;
  assign ram_b_7_0_enable = (_mystream_stream_oready && _mystream_b7_source_ram_renable && (_mystream_b7_source_sel == 40))? 1'd1 : 
                            ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  localparam _tmp_303 = 1;
  wire [_tmp_303-1:0] _tmp_304;
  assign _tmp_304 = _mystream_stream_oready && _mystream_b7_source_ram_renable && (_mystream_b7_source_sel == 40);
  reg [_tmp_303-1:0] __tmp_304_1;
  assign _mystream_b7_source_ram_rdata = (_mystream_b7_source_sel == 40)? ram_b_7_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_41;
  assign mystream_b7_data = __variable_wdata_41;
  reg [32-1:0] _mystream_b7_source_fsm_39;
  localparam _mystream_b7_source_fsm_39_init = 0;
  wire _set_flag_305;
  assign _set_flag_305 = th_comp == 56;
  assign ram_b_8_0_addr = (_mystream_stream_oready && _mystream_b8_source_ram_renable && (_mystream_b8_source_sel == 41))? _mystream_b8_source_ram_raddr : 
                          ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_addr_135 : 'hx;
  assign ram_b_8_0_enable = (_mystream_stream_oready && _mystream_b8_source_ram_renable && (_mystream_b8_source_sel == 41))? 1'd1 : 
                            ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  localparam _tmp_306 = 1;
  wire [_tmp_306-1:0] _tmp_307;
  assign _tmp_307 = _mystream_stream_oready && _mystream_b8_source_ram_renable && (_mystream_b8_source_sel == 41);
  reg [_tmp_306-1:0] __tmp_307_1;
  assign _mystream_b8_source_ram_rdata = (_mystream_b8_source_sel == 41)? ram_b_8_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_42;
  assign mystream_b8_data = __variable_wdata_42;
  reg [32-1:0] _mystream_b8_source_fsm_40;
  localparam _mystream_b8_source_fsm_40_init = 0;
  wire _set_flag_308;
  assign _set_flag_308 = th_comp == 57;
  assign ram_b_9_0_addr = (_mystream_stream_oready && _mystream_b9_source_ram_renable && (_mystream_b9_source_sel == 42))? _mystream_b9_source_ram_raddr : 
                          ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_addr_137 : 'hx;
  assign ram_b_9_0_enable = (_mystream_stream_oready && _mystream_b9_source_ram_renable && (_mystream_b9_source_sel == 42))? 1'd1 : 
                            ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  localparam _tmp_309 = 1;
  wire [_tmp_309-1:0] _tmp_310;
  assign _tmp_310 = _mystream_stream_oready && _mystream_b9_source_ram_renable && (_mystream_b9_source_sel == 42);
  reg [_tmp_309-1:0] __tmp_310_1;
  assign _mystream_b9_source_ram_rdata = (_mystream_b9_source_sel == 42)? ram_b_9_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_43;
  assign mystream_b9_data = __variable_wdata_43;
  reg [32-1:0] _mystream_b9_source_fsm_41;
  localparam _mystream_b9_source_fsm_41_init = 0;
  wire _set_flag_311;
  assign _set_flag_311 = th_comp == 58;
  assign ram_b_10_0_addr = (_mystream_stream_oready && _mystream_b10_source_ram_renable && (_mystream_b10_source_sel == 43))? _mystream_b10_source_ram_raddr : 
                           ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_addr_139 : 'hx;
  assign ram_b_10_0_enable = (_mystream_stream_oready && _mystream_b10_source_ram_renable && (_mystream_b10_source_sel == 43))? 1'd1 : 
                             ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  localparam _tmp_312 = 1;
  wire [_tmp_312-1:0] _tmp_313;
  assign _tmp_313 = _mystream_stream_oready && _mystream_b10_source_ram_renable && (_mystream_b10_source_sel == 43);
  reg [_tmp_312-1:0] __tmp_313_1;
  assign _mystream_b10_source_ram_rdata = (_mystream_b10_source_sel == 43)? ram_b_10_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_44;
  assign mystream_b10_data = __variable_wdata_44;
  reg [32-1:0] _mystream_b10_source_fsm_42;
  localparam _mystream_b10_source_fsm_42_init = 0;
  wire _set_flag_314;
  assign _set_flag_314 = th_comp == 59;
  assign ram_b_11_0_addr = (_mystream_stream_oready && _mystream_b11_source_ram_renable && (_mystream_b11_source_sel == 44))? _mystream_b11_source_ram_raddr : 
                           ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_addr_141 : 'hx;
  assign ram_b_11_0_enable = (_mystream_stream_oready && _mystream_b11_source_ram_renable && (_mystream_b11_source_sel == 44))? 1'd1 : 
                             ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  localparam _tmp_315 = 1;
  wire [_tmp_315-1:0] _tmp_316;
  assign _tmp_316 = _mystream_stream_oready && _mystream_b11_source_ram_renable && (_mystream_b11_source_sel == 44);
  reg [_tmp_315-1:0] __tmp_316_1;
  assign _mystream_b11_source_ram_rdata = (_mystream_b11_source_sel == 44)? ram_b_11_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_45;
  assign mystream_b11_data = __variable_wdata_45;
  reg [32-1:0] _mystream_b11_source_fsm_43;
  localparam _mystream_b11_source_fsm_43_init = 0;
  wire _set_flag_317;
  assign _set_flag_317 = th_comp == 60;
  assign ram_b_12_0_addr = (_mystream_stream_oready && _mystream_b12_source_ram_renable && (_mystream_b12_source_sel == 45))? _mystream_b12_source_ram_raddr : 
                           ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_addr_143 : 'hx;
  assign ram_b_12_0_enable = (_mystream_stream_oready && _mystream_b12_source_ram_renable && (_mystream_b12_source_sel == 45))? 1'd1 : 
                             ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  localparam _tmp_318 = 1;
  wire [_tmp_318-1:0] _tmp_319;
  assign _tmp_319 = _mystream_stream_oready && _mystream_b12_source_ram_renable && (_mystream_b12_source_sel == 45);
  reg [_tmp_318-1:0] __tmp_319_1;
  assign _mystream_b12_source_ram_rdata = (_mystream_b12_source_sel == 45)? ram_b_12_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_46;
  assign mystream_b12_data = __variable_wdata_46;
  reg [32-1:0] _mystream_b12_source_fsm_44;
  localparam _mystream_b12_source_fsm_44_init = 0;
  wire _set_flag_320;
  assign _set_flag_320 = th_comp == 61;
  assign ram_b_13_0_addr = (_mystream_stream_oready && _mystream_b13_source_ram_renable && (_mystream_b13_source_sel == 46))? _mystream_b13_source_ram_raddr : 
                           ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_addr_145 : 'hx;
  assign ram_b_13_0_enable = (_mystream_stream_oready && _mystream_b13_source_ram_renable && (_mystream_b13_source_sel == 46))? 1'd1 : 
                             ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  localparam _tmp_321 = 1;
  wire [_tmp_321-1:0] _tmp_322;
  assign _tmp_322 = _mystream_stream_oready && _mystream_b13_source_ram_renable && (_mystream_b13_source_sel == 46);
  reg [_tmp_321-1:0] __tmp_322_1;
  assign _mystream_b13_source_ram_rdata = (_mystream_b13_source_sel == 46)? ram_b_13_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_47;
  assign mystream_b13_data = __variable_wdata_47;
  reg [32-1:0] _mystream_b13_source_fsm_45;
  localparam _mystream_b13_source_fsm_45_init = 0;
  wire _set_flag_323;
  assign _set_flag_323 = th_comp == 62;
  assign ram_b_14_0_addr = (_mystream_stream_oready && _mystream_b14_source_ram_renable && (_mystream_b14_source_sel == 47))? _mystream_b14_source_ram_raddr : 
                           ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_addr_147 : 'hx;
  assign ram_b_14_0_enable = (_mystream_stream_oready && _mystream_b14_source_ram_renable && (_mystream_b14_source_sel == 47))? 1'd1 : 
                             ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  localparam _tmp_324 = 1;
  wire [_tmp_324-1:0] _tmp_325;
  assign _tmp_325 = _mystream_stream_oready && _mystream_b14_source_ram_renable && (_mystream_b14_source_sel == 47);
  reg [_tmp_324-1:0] __tmp_325_1;
  assign _mystream_b14_source_ram_rdata = (_mystream_b14_source_sel == 47)? ram_b_14_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_48;
  assign mystream_b14_data = __variable_wdata_48;
  reg [32-1:0] _mystream_b14_source_fsm_46;
  localparam _mystream_b14_source_fsm_46_init = 0;
  wire _set_flag_326;
  assign _set_flag_326 = th_comp == 63;
  assign ram_b_15_0_addr = (_mystream_stream_oready && _mystream_b15_source_ram_renable && (_mystream_b15_source_sel == 48))? _mystream_b15_source_ram_raddr : 
                           ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_addr_149 : 'hx;
  assign ram_b_15_0_enable = (_mystream_stream_oready && _mystream_b15_source_ram_renable && (_mystream_b15_source_sel == 48))? 1'd1 : 
                             ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  localparam _tmp_327 = 1;
  wire [_tmp_327-1:0] _tmp_328;
  assign _tmp_328 = _mystream_stream_oready && _mystream_b15_source_ram_renable && (_mystream_b15_source_sel == 48);
  reg [_tmp_327-1:0] __tmp_328_1;
  assign _mystream_b15_source_ram_rdata = (_mystream_b15_source_sel == 48)? ram_b_15_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_49;
  assign mystream_b15_data = __variable_wdata_49;
  reg [32-1:0] _mystream_b15_source_fsm_47;
  localparam _mystream_b15_source_fsm_47_init = 0;
  wire _set_flag_329;
  assign _set_flag_329 = th_comp == 64;
  assign ram_b_16_0_addr = (_mystream_stream_oready && _mystream_b16_source_ram_renable && (_mystream_b16_source_sel == 49))? _mystream_b16_source_ram_raddr : 
                           ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_addr_151 : 'hx;
  assign ram_b_16_0_enable = (_mystream_stream_oready && _mystream_b16_source_ram_renable && (_mystream_b16_source_sel == 49))? 1'd1 : 
                             ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  localparam _tmp_330 = 1;
  wire [_tmp_330-1:0] _tmp_331;
  assign _tmp_331 = _mystream_stream_oready && _mystream_b16_source_ram_renable && (_mystream_b16_source_sel == 49);
  reg [_tmp_330-1:0] __tmp_331_1;
  assign _mystream_b16_source_ram_rdata = (_mystream_b16_source_sel == 49)? ram_b_16_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_50;
  assign mystream_b16_data = __variable_wdata_50;
  reg [32-1:0] _mystream_b16_source_fsm_48;
  localparam _mystream_b16_source_fsm_48_init = 0;
  wire _set_flag_332;
  assign _set_flag_332 = th_comp == 65;
  assign ram_b_17_0_addr = (_mystream_stream_oready && _mystream_b17_source_ram_renable && (_mystream_b17_source_sel == 50))? _mystream_b17_source_ram_raddr : 
                           ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_addr_153 : 'hx;
  assign ram_b_17_0_enable = (_mystream_stream_oready && _mystream_b17_source_ram_renable && (_mystream_b17_source_sel == 50))? 1'd1 : 
                             ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  localparam _tmp_333 = 1;
  wire [_tmp_333-1:0] _tmp_334;
  assign _tmp_334 = _mystream_stream_oready && _mystream_b17_source_ram_renable && (_mystream_b17_source_sel == 50);
  reg [_tmp_333-1:0] __tmp_334_1;
  assign _mystream_b17_source_ram_rdata = (_mystream_b17_source_sel == 50)? ram_b_17_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_51;
  assign mystream_b17_data = __variable_wdata_51;
  reg [32-1:0] _mystream_b17_source_fsm_49;
  localparam _mystream_b17_source_fsm_49_init = 0;
  wire _set_flag_335;
  assign _set_flag_335 = th_comp == 66;
  assign ram_b_18_0_addr = (_mystream_stream_oready && _mystream_b18_source_ram_renable && (_mystream_b18_source_sel == 51))? _mystream_b18_source_ram_raddr : 
                           ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_addr_155 : 'hx;
  assign ram_b_18_0_enable = (_mystream_stream_oready && _mystream_b18_source_ram_renable && (_mystream_b18_source_sel == 51))? 1'd1 : 
                             ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  localparam _tmp_336 = 1;
  wire [_tmp_336-1:0] _tmp_337;
  assign _tmp_337 = _mystream_stream_oready && _mystream_b18_source_ram_renable && (_mystream_b18_source_sel == 51);
  reg [_tmp_336-1:0] __tmp_337_1;
  assign _mystream_b18_source_ram_rdata = (_mystream_b18_source_sel == 51)? ram_b_18_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_52;
  assign mystream_b18_data = __variable_wdata_52;
  reg [32-1:0] _mystream_b18_source_fsm_50;
  localparam _mystream_b18_source_fsm_50_init = 0;
  wire _set_flag_338;
  assign _set_flag_338 = th_comp == 67;
  assign ram_b_19_0_addr = (_mystream_stream_oready && _mystream_b19_source_ram_renable && (_mystream_b19_source_sel == 52))? _mystream_b19_source_ram_raddr : 
                           ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_addr_157 : 'hx;
  assign ram_b_19_0_enable = (_mystream_stream_oready && _mystream_b19_source_ram_renable && (_mystream_b19_source_sel == 52))? 1'd1 : 
                             ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  localparam _tmp_339 = 1;
  wire [_tmp_339-1:0] _tmp_340;
  assign _tmp_340 = _mystream_stream_oready && _mystream_b19_source_ram_renable && (_mystream_b19_source_sel == 52);
  reg [_tmp_339-1:0] __tmp_340_1;
  assign _mystream_b19_source_ram_rdata = (_mystream_b19_source_sel == 52)? ram_b_19_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_53;
  assign mystream_b19_data = __variable_wdata_53;
  reg [32-1:0] _mystream_b19_source_fsm_51;
  localparam _mystream_b19_source_fsm_51_init = 0;
  wire _set_flag_341;
  assign _set_flag_341 = th_comp == 68;
  assign ram_b_20_0_addr = (_mystream_stream_oready && _mystream_b20_source_ram_renable && (_mystream_b20_source_sel == 53))? _mystream_b20_source_ram_raddr : 
                           ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_addr_159 : 'hx;
  assign ram_b_20_0_enable = (_mystream_stream_oready && _mystream_b20_source_ram_renable && (_mystream_b20_source_sel == 53))? 1'd1 : 
                             ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  localparam _tmp_342 = 1;
  wire [_tmp_342-1:0] _tmp_343;
  assign _tmp_343 = _mystream_stream_oready && _mystream_b20_source_ram_renable && (_mystream_b20_source_sel == 53);
  reg [_tmp_342-1:0] __tmp_343_1;
  assign _mystream_b20_source_ram_rdata = (_mystream_b20_source_sel == 53)? ram_b_20_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_54;
  assign mystream_b20_data = __variable_wdata_54;
  reg [32-1:0] _mystream_b20_source_fsm_52;
  localparam _mystream_b20_source_fsm_52_init = 0;
  wire _set_flag_344;
  assign _set_flag_344 = th_comp == 69;
  assign ram_b_21_0_addr = (_mystream_stream_oready && _mystream_b21_source_ram_renable && (_mystream_b21_source_sel == 54))? _mystream_b21_source_ram_raddr : 
                           ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_addr_161 : 'hx;
  assign ram_b_21_0_enable = (_mystream_stream_oready && _mystream_b21_source_ram_renable && (_mystream_b21_source_sel == 54))? 1'd1 : 
                             ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  localparam _tmp_345 = 1;
  wire [_tmp_345-1:0] _tmp_346;
  assign _tmp_346 = _mystream_stream_oready && _mystream_b21_source_ram_renable && (_mystream_b21_source_sel == 54);
  reg [_tmp_345-1:0] __tmp_346_1;
  assign _mystream_b21_source_ram_rdata = (_mystream_b21_source_sel == 54)? ram_b_21_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_55;
  assign mystream_b21_data = __variable_wdata_55;
  reg [32-1:0] _mystream_b21_source_fsm_53;
  localparam _mystream_b21_source_fsm_53_init = 0;
  wire _set_flag_347;
  assign _set_flag_347 = th_comp == 70;
  assign ram_b_22_0_addr = (_mystream_stream_oready && _mystream_b22_source_ram_renable && (_mystream_b22_source_sel == 55))? _mystream_b22_source_ram_raddr : 
                           ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_addr_163 : 'hx;
  assign ram_b_22_0_enable = (_mystream_stream_oready && _mystream_b22_source_ram_renable && (_mystream_b22_source_sel == 55))? 1'd1 : 
                             ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  localparam _tmp_348 = 1;
  wire [_tmp_348-1:0] _tmp_349;
  assign _tmp_349 = _mystream_stream_oready && _mystream_b22_source_ram_renable && (_mystream_b22_source_sel == 55);
  reg [_tmp_348-1:0] __tmp_349_1;
  assign _mystream_b22_source_ram_rdata = (_mystream_b22_source_sel == 55)? ram_b_22_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_56;
  assign mystream_b22_data = __variable_wdata_56;
  reg [32-1:0] _mystream_b22_source_fsm_54;
  localparam _mystream_b22_source_fsm_54_init = 0;
  wire _set_flag_350;
  assign _set_flag_350 = th_comp == 71;
  assign ram_b_23_0_addr = (_mystream_stream_oready && _mystream_b23_source_ram_renable && (_mystream_b23_source_sel == 56))? _mystream_b23_source_ram_raddr : 
                           ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_addr_165 : 'hx;
  assign ram_b_23_0_enable = (_mystream_stream_oready && _mystream_b23_source_ram_renable && (_mystream_b23_source_sel == 56))? 1'd1 : 
                             ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  localparam _tmp_351 = 1;
  wire [_tmp_351-1:0] _tmp_352;
  assign _tmp_352 = _mystream_stream_oready && _mystream_b23_source_ram_renable && (_mystream_b23_source_sel == 56);
  reg [_tmp_351-1:0] __tmp_352_1;
  assign _mystream_b23_source_ram_rdata = (_mystream_b23_source_sel == 56)? ram_b_23_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_57;
  assign mystream_b23_data = __variable_wdata_57;
  reg [32-1:0] _mystream_b23_source_fsm_55;
  localparam _mystream_b23_source_fsm_55_init = 0;
  wire _set_flag_353;
  assign _set_flag_353 = th_comp == 72;
  assign ram_b_24_0_addr = (_mystream_stream_oready && _mystream_b24_source_ram_renable && (_mystream_b24_source_sel == 57))? _mystream_b24_source_ram_raddr : 
                           ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_addr_167 : 'hx;
  assign ram_b_24_0_enable = (_mystream_stream_oready && _mystream_b24_source_ram_renable && (_mystream_b24_source_sel == 57))? 1'd1 : 
                             ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  localparam _tmp_354 = 1;
  wire [_tmp_354-1:0] _tmp_355;
  assign _tmp_355 = _mystream_stream_oready && _mystream_b24_source_ram_renable && (_mystream_b24_source_sel == 57);
  reg [_tmp_354-1:0] __tmp_355_1;
  assign _mystream_b24_source_ram_rdata = (_mystream_b24_source_sel == 57)? ram_b_24_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_58;
  assign mystream_b24_data = __variable_wdata_58;
  reg [32-1:0] _mystream_b24_source_fsm_56;
  localparam _mystream_b24_source_fsm_56_init = 0;
  wire _set_flag_356;
  assign _set_flag_356 = th_comp == 73;
  assign ram_b_25_0_addr = (_mystream_stream_oready && _mystream_b25_source_ram_renable && (_mystream_b25_source_sel == 58))? _mystream_b25_source_ram_raddr : 
                           ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_addr_169 : 'hx;
  assign ram_b_25_0_enable = (_mystream_stream_oready && _mystream_b25_source_ram_renable && (_mystream_b25_source_sel == 58))? 1'd1 : 
                             ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  localparam _tmp_357 = 1;
  wire [_tmp_357-1:0] _tmp_358;
  assign _tmp_358 = _mystream_stream_oready && _mystream_b25_source_ram_renable && (_mystream_b25_source_sel == 58);
  reg [_tmp_357-1:0] __tmp_358_1;
  assign _mystream_b25_source_ram_rdata = (_mystream_b25_source_sel == 58)? ram_b_25_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_59;
  assign mystream_b25_data = __variable_wdata_59;
  reg [32-1:0] _mystream_b25_source_fsm_57;
  localparam _mystream_b25_source_fsm_57_init = 0;
  wire _set_flag_359;
  assign _set_flag_359 = th_comp == 74;
  assign ram_b_26_0_addr = (_mystream_stream_oready && _mystream_b26_source_ram_renable && (_mystream_b26_source_sel == 59))? _mystream_b26_source_ram_raddr : 
                           ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_addr_171 : 'hx;
  assign ram_b_26_0_enable = (_mystream_stream_oready && _mystream_b26_source_ram_renable && (_mystream_b26_source_sel == 59))? 1'd1 : 
                             ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  localparam _tmp_360 = 1;
  wire [_tmp_360-1:0] _tmp_361;
  assign _tmp_361 = _mystream_stream_oready && _mystream_b26_source_ram_renable && (_mystream_b26_source_sel == 59);
  reg [_tmp_360-1:0] __tmp_361_1;
  assign _mystream_b26_source_ram_rdata = (_mystream_b26_source_sel == 59)? ram_b_26_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_60;
  assign mystream_b26_data = __variable_wdata_60;
  reg [32-1:0] _mystream_b26_source_fsm_58;
  localparam _mystream_b26_source_fsm_58_init = 0;
  wire _set_flag_362;
  assign _set_flag_362 = th_comp == 75;
  assign ram_b_27_0_addr = (_mystream_stream_oready && _mystream_b27_source_ram_renable && (_mystream_b27_source_sel == 60))? _mystream_b27_source_ram_raddr : 
                           ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_addr_173 : 'hx;
  assign ram_b_27_0_enable = (_mystream_stream_oready && _mystream_b27_source_ram_renable && (_mystream_b27_source_sel == 60))? 1'd1 : 
                             ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  localparam _tmp_363 = 1;
  wire [_tmp_363-1:0] _tmp_364;
  assign _tmp_364 = _mystream_stream_oready && _mystream_b27_source_ram_renable && (_mystream_b27_source_sel == 60);
  reg [_tmp_363-1:0] __tmp_364_1;
  assign _mystream_b27_source_ram_rdata = (_mystream_b27_source_sel == 60)? ram_b_27_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_61;
  assign mystream_b27_data = __variable_wdata_61;
  reg [32-1:0] _mystream_b27_source_fsm_59;
  localparam _mystream_b27_source_fsm_59_init = 0;
  wire _set_flag_365;
  assign _set_flag_365 = th_comp == 76;
  assign ram_b_28_0_addr = (_mystream_stream_oready && _mystream_b28_source_ram_renable && (_mystream_b28_source_sel == 61))? _mystream_b28_source_ram_raddr : 
                           ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_addr_175 : 'hx;
  assign ram_b_28_0_enable = (_mystream_stream_oready && _mystream_b28_source_ram_renable && (_mystream_b28_source_sel == 61))? 1'd1 : 
                             ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  localparam _tmp_366 = 1;
  wire [_tmp_366-1:0] _tmp_367;
  assign _tmp_367 = _mystream_stream_oready && _mystream_b28_source_ram_renable && (_mystream_b28_source_sel == 61);
  reg [_tmp_366-1:0] __tmp_367_1;
  assign _mystream_b28_source_ram_rdata = (_mystream_b28_source_sel == 61)? ram_b_28_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_62;
  assign mystream_b28_data = __variable_wdata_62;
  reg [32-1:0] _mystream_b28_source_fsm_60;
  localparam _mystream_b28_source_fsm_60_init = 0;
  wire _set_flag_368;
  assign _set_flag_368 = th_comp == 77;
  assign ram_b_29_0_addr = (_mystream_stream_oready && _mystream_b29_source_ram_renable && (_mystream_b29_source_sel == 62))? _mystream_b29_source_ram_raddr : 
                           ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_addr_177 : 'hx;
  assign ram_b_29_0_enable = (_mystream_stream_oready && _mystream_b29_source_ram_renable && (_mystream_b29_source_sel == 62))? 1'd1 : 
                             ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  localparam _tmp_369 = 1;
  wire [_tmp_369-1:0] _tmp_370;
  assign _tmp_370 = _mystream_stream_oready && _mystream_b29_source_ram_renable && (_mystream_b29_source_sel == 62);
  reg [_tmp_369-1:0] __tmp_370_1;
  assign _mystream_b29_source_ram_rdata = (_mystream_b29_source_sel == 62)? ram_b_29_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_63;
  assign mystream_b29_data = __variable_wdata_63;
  reg [32-1:0] _mystream_b29_source_fsm_61;
  localparam _mystream_b29_source_fsm_61_init = 0;
  wire _set_flag_371;
  assign _set_flag_371 = th_comp == 78;
  assign ram_b_30_0_addr = (_mystream_stream_oready && _mystream_b30_source_ram_renable && (_mystream_b30_source_sel == 63))? _mystream_b30_source_ram_raddr : 
                           ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_addr_179 : 'hx;
  assign ram_b_30_0_enable = (_mystream_stream_oready && _mystream_b30_source_ram_renable && (_mystream_b30_source_sel == 63))? 1'd1 : 
                             ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  localparam _tmp_372 = 1;
  wire [_tmp_372-1:0] _tmp_373;
  assign _tmp_373 = _mystream_stream_oready && _mystream_b30_source_ram_renable && (_mystream_b30_source_sel == 63);
  reg [_tmp_372-1:0] __tmp_373_1;
  assign _mystream_b30_source_ram_rdata = (_mystream_b30_source_sel == 63)? ram_b_30_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_64;
  assign mystream_b30_data = __variable_wdata_64;
  reg [32-1:0] _mystream_b30_source_fsm_62;
  localparam _mystream_b30_source_fsm_62_init = 0;
  wire _set_flag_374;
  assign _set_flag_374 = th_comp == 79;
  assign ram_b_31_0_addr = (_mystream_stream_oready && _mystream_b31_source_ram_renable && (_mystream_b31_source_sel == 64))? _mystream_b31_source_ram_raddr : 
                           ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? write_burst_packed_ram_addr_181 : 'hx;
  assign ram_b_31_0_enable = (_mystream_stream_oready && _mystream_b31_source_ram_renable && (_mystream_b31_source_sel == 64))? 1'd1 : 
                             ((write_burst_packed_fsm_1 == 1) && _myaxi_read_narrow_wvalid_113)? 1'd1 : 0;
  localparam _tmp_375 = 1;
  wire [_tmp_375-1:0] _tmp_376;
  assign _tmp_376 = _mystream_stream_oready && _mystream_b31_source_ram_renable && (_mystream_b31_source_sel == 64);
  reg [_tmp_375-1:0] __tmp_376_1;
  assign _mystream_b31_source_ram_rdata = (_mystream_b31_source_sel == 64)? ram_b_31_0_rdata : 'hx;
  reg signed [32-1:0] __variable_wdata_65;
  assign mystream_b31_data = __variable_wdata_65;
  reg [32-1:0] _mystream_b31_source_fsm_63;
  localparam _mystream_b31_source_fsm_63_init = 0;
  wire _set_flag_377;
  assign _set_flag_377 = th_comp == 82;
  reg _tmp_378;
  reg _tmp_379;
  reg _tmp_380;
  reg _tmp_381;
  reg _tmp_382;
  reg _tmp_383;
  reg signed [32-1:0] _tmp_384;
  reg signed [32-1:0] _tmp_385;
  reg signed [32-1:0] _tmp_386;
  reg signed [32-1:0] _tmp_387;
  reg signed [32-1:0] _tmp_388;
  reg signed [32-1:0] _tmp_389;
  localparam _tmp_390 = 34;
  wire [_tmp_390-1:0] _tmp_391;
  assign _tmp_391 = _th_comp_size_3 + 32 - 1 >>> 5;
  reg [_tmp_390-1:0] _tmp_392;
  reg [_tmp_390-1:0] _tmp_393;
  reg [_tmp_390-1:0] _tmp_394;
  reg [_tmp_390-1:0] _tmp_395;
  reg [_tmp_390-1:0] _tmp_396;
  reg [_tmp_390-1:0] _tmp_397;
  reg [32-1:0] _mystream_sum_vec0_sink_fsm_64;
  localparam _mystream_sum_vec0_sink_fsm_64_init = 0;
  wire _set_flag_398;
  assign _set_flag_398 = th_comp == 82;
  reg _tmp_399;
  reg _tmp_400;
  reg _tmp_401;
  reg _tmp_402;
  reg _tmp_403;
  reg _tmp_404;
  reg signed [32-1:0] _tmp_405;
  reg signed [32-1:0] _tmp_406;
  reg signed [32-1:0] _tmp_407;
  reg signed [32-1:0] _tmp_408;
  reg signed [32-1:0] _tmp_409;
  reg signed [32-1:0] _tmp_410;
  localparam _tmp_411 = 34;
  wire [_tmp_411-1:0] _tmp_412;
  assign _tmp_412 = _th_comp_size_3 + 32 - 1 >>> 5;
  reg [_tmp_411-1:0] _tmp_413;
  reg [_tmp_411-1:0] _tmp_414;
  reg [_tmp_411-1:0] _tmp_415;
  reg [_tmp_411-1:0] _tmp_416;
  reg [_tmp_411-1:0] _tmp_417;
  reg [_tmp_411-1:0] _tmp_418;
  reg [32-1:0] _mystream_sum_vec1_sink_fsm_65;
  localparam _mystream_sum_vec1_sink_fsm_65_init = 0;
  wire _set_flag_419;
  assign _set_flag_419 = th_comp == 82;
  reg _tmp_420;
  reg _tmp_421;
  reg _tmp_422;
  reg _tmp_423;
  reg _tmp_424;
  reg _tmp_425;
  reg signed [32-1:0] _tmp_426;
  reg signed [32-1:0] _tmp_427;
  reg signed [32-1:0] _tmp_428;
  reg signed [32-1:0] _tmp_429;
  reg signed [32-1:0] _tmp_430;
  reg signed [32-1:0] _tmp_431;
  localparam _tmp_432 = 34;
  wire [_tmp_432-1:0] _tmp_433;
  assign _tmp_433 = _th_comp_size_3 + 32 - 1 >>> 5;
  reg [_tmp_432-1:0] _tmp_434;
  reg [_tmp_432-1:0] _tmp_435;
  reg [_tmp_432-1:0] _tmp_436;
  reg [_tmp_432-1:0] _tmp_437;
  reg [_tmp_432-1:0] _tmp_438;
  reg [_tmp_432-1:0] _tmp_439;
  reg [32-1:0] _mystream_sum_vec2_sink_fsm_66;
  localparam _mystream_sum_vec2_sink_fsm_66_init = 0;
  wire _set_flag_440;
  assign _set_flag_440 = th_comp == 82;
  reg _tmp_441;
  reg _tmp_442;
  reg _tmp_443;
  reg _tmp_444;
  reg _tmp_445;
  reg _tmp_446;
  reg signed [32-1:0] _tmp_447;
  reg signed [32-1:0] _tmp_448;
  reg signed [32-1:0] _tmp_449;
  reg signed [32-1:0] _tmp_450;
  reg signed [32-1:0] _tmp_451;
  reg signed [32-1:0] _tmp_452;
  localparam _tmp_453 = 34;
  wire [_tmp_453-1:0] _tmp_454;
  assign _tmp_454 = _th_comp_size_3 + 32 - 1 >>> 5;
  reg [_tmp_453-1:0] _tmp_455;
  reg [_tmp_453-1:0] _tmp_456;
  reg [_tmp_453-1:0] _tmp_457;
  reg [_tmp_453-1:0] _tmp_458;
  reg [_tmp_453-1:0] _tmp_459;
  reg [_tmp_453-1:0] _tmp_460;
  reg [32-1:0] _mystream_sum_vec3_sink_fsm_67;
  localparam _mystream_sum_vec3_sink_fsm_67_init = 0;
  wire _set_flag_461;
  assign _set_flag_461 = th_comp == 82;
  reg _tmp_462;
  reg _tmp_463;
  reg _tmp_464;
  reg _tmp_465;
  reg _tmp_466;
  reg _tmp_467;
  reg signed [32-1:0] _tmp_468;
  reg signed [32-1:0] _tmp_469;
  reg signed [32-1:0] _tmp_470;
  reg signed [32-1:0] _tmp_471;
  reg signed [32-1:0] _tmp_472;
  reg signed [32-1:0] _tmp_473;
  localparam _tmp_474 = 34;
  wire [_tmp_474-1:0] _tmp_475;
  assign _tmp_475 = _th_comp_size_3 + 32 - 1 >>> 5;
  reg [_tmp_474-1:0] _tmp_476;
  reg [_tmp_474-1:0] _tmp_477;
  reg [_tmp_474-1:0] _tmp_478;
  reg [_tmp_474-1:0] _tmp_479;
  reg [_tmp_474-1:0] _tmp_480;
  reg [_tmp_474-1:0] _tmp_481;
  reg [32-1:0] _mystream_sum_vec4_sink_fsm_68;
  localparam _mystream_sum_vec4_sink_fsm_68_init = 0;
  wire _set_flag_482;
  assign _set_flag_482 = th_comp == 82;
  reg _tmp_483;
  reg _tmp_484;
  reg _tmp_485;
  reg _tmp_486;
  reg _tmp_487;
  reg _tmp_488;
  reg signed [32-1:0] _tmp_489;
  reg signed [32-1:0] _tmp_490;
  reg signed [32-1:0] _tmp_491;
  reg signed [32-1:0] _tmp_492;
  reg signed [32-1:0] _tmp_493;
  reg signed [32-1:0] _tmp_494;
  localparam _tmp_495 = 34;
  wire [_tmp_495-1:0] _tmp_496;
  assign _tmp_496 = _th_comp_size_3 + 32 - 1 >>> 5;
  reg [_tmp_495-1:0] _tmp_497;
  reg [_tmp_495-1:0] _tmp_498;
  reg [_tmp_495-1:0] _tmp_499;
  reg [_tmp_495-1:0] _tmp_500;
  reg [_tmp_495-1:0] _tmp_501;
  reg [_tmp_495-1:0] _tmp_502;
  reg [32-1:0] _mystream_sum_vec5_sink_fsm_69;
  localparam _mystream_sum_vec5_sink_fsm_69_init = 0;
  wire _set_flag_503;
  assign _set_flag_503 = th_comp == 82;
  reg _tmp_504;
  reg _tmp_505;
  reg _tmp_506;
  reg _tmp_507;
  reg _tmp_508;
  reg _tmp_509;
  reg signed [32-1:0] _tmp_510;
  reg signed [32-1:0] _tmp_511;
  reg signed [32-1:0] _tmp_512;
  reg signed [32-1:0] _tmp_513;
  reg signed [32-1:0] _tmp_514;
  reg signed [32-1:0] _tmp_515;
  localparam _tmp_516 = 34;
  wire [_tmp_516-1:0] _tmp_517;
  assign _tmp_517 = _th_comp_size_3 + 32 - 1 >>> 5;
  reg [_tmp_516-1:0] _tmp_518;
  reg [_tmp_516-1:0] _tmp_519;
  reg [_tmp_516-1:0] _tmp_520;
  reg [_tmp_516-1:0] _tmp_521;
  reg [_tmp_516-1:0] _tmp_522;
  reg [_tmp_516-1:0] _tmp_523;
  reg [32-1:0] _mystream_sum_vec6_sink_fsm_70;
  localparam _mystream_sum_vec6_sink_fsm_70_init = 0;
  wire _set_flag_524;
  assign _set_flag_524 = th_comp == 82;
  reg _tmp_525;
  reg _tmp_526;
  reg _tmp_527;
  reg _tmp_528;
  reg _tmp_529;
  reg _tmp_530;
  reg signed [32-1:0] _tmp_531;
  reg signed [32-1:0] _tmp_532;
  reg signed [32-1:0] _tmp_533;
  reg signed [32-1:0] _tmp_534;
  reg signed [32-1:0] _tmp_535;
  reg signed [32-1:0] _tmp_536;
  localparam _tmp_537 = 34;
  wire [_tmp_537-1:0] _tmp_538;
  assign _tmp_538 = _th_comp_size_3 + 32 - 1 >>> 5;
  reg [_tmp_537-1:0] _tmp_539;
  reg [_tmp_537-1:0] _tmp_540;
  reg [_tmp_537-1:0] _tmp_541;
  reg [_tmp_537-1:0] _tmp_542;
  reg [_tmp_537-1:0] _tmp_543;
  reg [_tmp_537-1:0] _tmp_544;
  reg [32-1:0] _mystream_sum_vec7_sink_fsm_71;
  localparam _mystream_sum_vec7_sink_fsm_71_init = 0;
  wire _set_flag_545;
  assign _set_flag_545 = th_comp == 82;
  reg _tmp_546;
  reg _tmp_547;
  reg _tmp_548;
  reg _tmp_549;
  reg _tmp_550;
  reg _tmp_551;
  reg signed [32-1:0] _tmp_552;
  reg signed [32-1:0] _tmp_553;
  reg signed [32-1:0] _tmp_554;
  reg signed [32-1:0] _tmp_555;
  reg signed [32-1:0] _tmp_556;
  reg signed [32-1:0] _tmp_557;
  localparam _tmp_558 = 34;
  wire [_tmp_558-1:0] _tmp_559;
  assign _tmp_559 = _th_comp_size_3 + 32 - 1 >>> 5;
  reg [_tmp_558-1:0] _tmp_560;
  reg [_tmp_558-1:0] _tmp_561;
  reg [_tmp_558-1:0] _tmp_562;
  reg [_tmp_558-1:0] _tmp_563;
  reg [_tmp_558-1:0] _tmp_564;
  reg [_tmp_558-1:0] _tmp_565;
  reg [32-1:0] _mystream_sum_vec8_sink_fsm_72;
  localparam _mystream_sum_vec8_sink_fsm_72_init = 0;
  wire _set_flag_566;
  assign _set_flag_566 = th_comp == 82;
  reg _tmp_567;
  reg _tmp_568;
  reg _tmp_569;
  reg _tmp_570;
  reg _tmp_571;
  reg _tmp_572;
  reg signed [32-1:0] _tmp_573;
  reg signed [32-1:0] _tmp_574;
  reg signed [32-1:0] _tmp_575;
  reg signed [32-1:0] _tmp_576;
  reg signed [32-1:0] _tmp_577;
  reg signed [32-1:0] _tmp_578;
  localparam _tmp_579 = 34;
  wire [_tmp_579-1:0] _tmp_580;
  assign _tmp_580 = _th_comp_size_3 + 32 - 1 >>> 5;
  reg [_tmp_579-1:0] _tmp_581;
  reg [_tmp_579-1:0] _tmp_582;
  reg [_tmp_579-1:0] _tmp_583;
  reg [_tmp_579-1:0] _tmp_584;
  reg [_tmp_579-1:0] _tmp_585;
  reg [_tmp_579-1:0] _tmp_586;
  reg [32-1:0] _mystream_sum_vec9_sink_fsm_73;
  localparam _mystream_sum_vec9_sink_fsm_73_init = 0;
  wire _set_flag_587;
  assign _set_flag_587 = th_comp == 82;
  reg _tmp_588;
  reg _tmp_589;
  reg _tmp_590;
  reg _tmp_591;
  reg _tmp_592;
  reg _tmp_593;
  reg signed [32-1:0] _tmp_594;
  reg signed [32-1:0] _tmp_595;
  reg signed [32-1:0] _tmp_596;
  reg signed [32-1:0] _tmp_597;
  reg signed [32-1:0] _tmp_598;
  reg signed [32-1:0] _tmp_599;
  localparam _tmp_600 = 34;
  wire [_tmp_600-1:0] _tmp_601;
  assign _tmp_601 = _th_comp_size_3 + 32 - 1 >>> 5;
  reg [_tmp_600-1:0] _tmp_602;
  reg [_tmp_600-1:0] _tmp_603;
  reg [_tmp_600-1:0] _tmp_604;
  reg [_tmp_600-1:0] _tmp_605;
  reg [_tmp_600-1:0] _tmp_606;
  reg [_tmp_600-1:0] _tmp_607;
  reg [32-1:0] _mystream_sum_vec10_sink_fsm_74;
  localparam _mystream_sum_vec10_sink_fsm_74_init = 0;
  wire _set_flag_608;
  assign _set_flag_608 = th_comp == 82;
  reg _tmp_609;
  reg _tmp_610;
  reg _tmp_611;
  reg _tmp_612;
  reg _tmp_613;
  reg _tmp_614;
  reg signed [32-1:0] _tmp_615;
  reg signed [32-1:0] _tmp_616;
  reg signed [32-1:0] _tmp_617;
  reg signed [32-1:0] _tmp_618;
  reg signed [32-1:0] _tmp_619;
  reg signed [32-1:0] _tmp_620;
  localparam _tmp_621 = 34;
  wire [_tmp_621-1:0] _tmp_622;
  assign _tmp_622 = _th_comp_size_3 + 32 - 1 >>> 5;
  reg [_tmp_621-1:0] _tmp_623;
  reg [_tmp_621-1:0] _tmp_624;
  reg [_tmp_621-1:0] _tmp_625;
  reg [_tmp_621-1:0] _tmp_626;
  reg [_tmp_621-1:0] _tmp_627;
  reg [_tmp_621-1:0] _tmp_628;
  reg [32-1:0] _mystream_sum_vec11_sink_fsm_75;
  localparam _mystream_sum_vec11_sink_fsm_75_init = 0;
  wire _set_flag_629;
  assign _set_flag_629 = th_comp == 82;
  reg _tmp_630;
  reg _tmp_631;
  reg _tmp_632;
  reg _tmp_633;
  reg _tmp_634;
  reg _tmp_635;
  reg signed [32-1:0] _tmp_636;
  reg signed [32-1:0] _tmp_637;
  reg signed [32-1:0] _tmp_638;
  reg signed [32-1:0] _tmp_639;
  reg signed [32-1:0] _tmp_640;
  reg signed [32-1:0] _tmp_641;
  localparam _tmp_642 = 34;
  wire [_tmp_642-1:0] _tmp_643;
  assign _tmp_643 = _th_comp_size_3 + 32 - 1 >>> 5;
  reg [_tmp_642-1:0] _tmp_644;
  reg [_tmp_642-1:0] _tmp_645;
  reg [_tmp_642-1:0] _tmp_646;
  reg [_tmp_642-1:0] _tmp_647;
  reg [_tmp_642-1:0] _tmp_648;
  reg [_tmp_642-1:0] _tmp_649;
  reg [32-1:0] _mystream_sum_vec12_sink_fsm_76;
  localparam _mystream_sum_vec12_sink_fsm_76_init = 0;
  wire _set_flag_650;
  assign _set_flag_650 = th_comp == 82;
  reg _tmp_651;
  reg _tmp_652;
  reg _tmp_653;
  reg _tmp_654;
  reg _tmp_655;
  reg _tmp_656;
  reg signed [32-1:0] _tmp_657;
  reg signed [32-1:0] _tmp_658;
  reg signed [32-1:0] _tmp_659;
  reg signed [32-1:0] _tmp_660;
  reg signed [32-1:0] _tmp_661;
  reg signed [32-1:0] _tmp_662;
  localparam _tmp_663 = 34;
  wire [_tmp_663-1:0] _tmp_664;
  assign _tmp_664 = _th_comp_size_3 + 32 - 1 >>> 5;
  reg [_tmp_663-1:0] _tmp_665;
  reg [_tmp_663-1:0] _tmp_666;
  reg [_tmp_663-1:0] _tmp_667;
  reg [_tmp_663-1:0] _tmp_668;
  reg [_tmp_663-1:0] _tmp_669;
  reg [_tmp_663-1:0] _tmp_670;
  reg [32-1:0] _mystream_sum_vec13_sink_fsm_77;
  localparam _mystream_sum_vec13_sink_fsm_77_init = 0;
  wire _set_flag_671;
  assign _set_flag_671 = th_comp == 82;
  reg _tmp_672;
  reg _tmp_673;
  reg _tmp_674;
  reg _tmp_675;
  reg _tmp_676;
  reg _tmp_677;
  reg signed [32-1:0] _tmp_678;
  reg signed [32-1:0] _tmp_679;
  reg signed [32-1:0] _tmp_680;
  reg signed [32-1:0] _tmp_681;
  reg signed [32-1:0] _tmp_682;
  reg signed [32-1:0] _tmp_683;
  localparam _tmp_684 = 34;
  wire [_tmp_684-1:0] _tmp_685;
  assign _tmp_685 = _th_comp_size_3 + 32 - 1 >>> 5;
  reg [_tmp_684-1:0] _tmp_686;
  reg [_tmp_684-1:0] _tmp_687;
  reg [_tmp_684-1:0] _tmp_688;
  reg [_tmp_684-1:0] _tmp_689;
  reg [_tmp_684-1:0] _tmp_690;
  reg [_tmp_684-1:0] _tmp_691;
  reg [32-1:0] _mystream_sum_vec14_sink_fsm_78;
  localparam _mystream_sum_vec14_sink_fsm_78_init = 0;
  wire _set_flag_692;
  assign _set_flag_692 = th_comp == 82;
  reg _tmp_693;
  reg _tmp_694;
  reg _tmp_695;
  reg _tmp_696;
  reg _tmp_697;
  reg _tmp_698;
  reg signed [32-1:0] _tmp_699;
  reg signed [32-1:0] _tmp_700;
  reg signed [32-1:0] _tmp_701;
  reg signed [32-1:0] _tmp_702;
  reg signed [32-1:0] _tmp_703;
  reg signed [32-1:0] _tmp_704;
  localparam _tmp_705 = 34;
  wire [_tmp_705-1:0] _tmp_706;
  assign _tmp_706 = _th_comp_size_3 + 32 - 1 >>> 5;
  reg [_tmp_705-1:0] _tmp_707;
  reg [_tmp_705-1:0] _tmp_708;
  reg [_tmp_705-1:0] _tmp_709;
  reg [_tmp_705-1:0] _tmp_710;
  reg [_tmp_705-1:0] _tmp_711;
  reg [_tmp_705-1:0] _tmp_712;
  reg [32-1:0] _mystream_sum_vec15_sink_fsm_79;
  localparam _mystream_sum_vec15_sink_fsm_79_init = 0;
  wire _set_flag_713;
  assign _set_flag_713 = th_comp == 82;
  reg _tmp_714;
  reg _tmp_715;
  reg _tmp_716;
  reg _tmp_717;
  reg _tmp_718;
  reg _tmp_719;
  reg signed [32-1:0] _tmp_720;
  reg signed [32-1:0] _tmp_721;
  reg signed [32-1:0] _tmp_722;
  reg signed [32-1:0] _tmp_723;
  reg signed [32-1:0] _tmp_724;
  reg signed [32-1:0] _tmp_725;
  localparam _tmp_726 = 34;
  wire [_tmp_726-1:0] _tmp_727;
  assign _tmp_727 = _th_comp_size_3 + 32 - 1 >>> 5;
  reg [_tmp_726-1:0] _tmp_728;
  reg [_tmp_726-1:0] _tmp_729;
  reg [_tmp_726-1:0] _tmp_730;
  reg [_tmp_726-1:0] _tmp_731;
  reg [_tmp_726-1:0] _tmp_732;
  reg [_tmp_726-1:0] _tmp_733;
  reg [32-1:0] _mystream_sum_vec16_sink_fsm_80;
  localparam _mystream_sum_vec16_sink_fsm_80_init = 0;
  wire _set_flag_734;
  assign _set_flag_734 = th_comp == 82;
  reg _tmp_735;
  reg _tmp_736;
  reg _tmp_737;
  reg _tmp_738;
  reg _tmp_739;
  reg _tmp_740;
  reg signed [32-1:0] _tmp_741;
  reg signed [32-1:0] _tmp_742;
  reg signed [32-1:0] _tmp_743;
  reg signed [32-1:0] _tmp_744;
  reg signed [32-1:0] _tmp_745;
  reg signed [32-1:0] _tmp_746;
  localparam _tmp_747 = 34;
  wire [_tmp_747-1:0] _tmp_748;
  assign _tmp_748 = _th_comp_size_3 + 32 - 1 >>> 5;
  reg [_tmp_747-1:0] _tmp_749;
  reg [_tmp_747-1:0] _tmp_750;
  reg [_tmp_747-1:0] _tmp_751;
  reg [_tmp_747-1:0] _tmp_752;
  reg [_tmp_747-1:0] _tmp_753;
  reg [_tmp_747-1:0] _tmp_754;
  reg [32-1:0] _mystream_sum_vec17_sink_fsm_81;
  localparam _mystream_sum_vec17_sink_fsm_81_init = 0;
  wire _set_flag_755;
  assign _set_flag_755 = th_comp == 82;
  reg _tmp_756;
  reg _tmp_757;
  reg _tmp_758;
  reg _tmp_759;
  reg _tmp_760;
  reg _tmp_761;
  reg signed [32-1:0] _tmp_762;
  reg signed [32-1:0] _tmp_763;
  reg signed [32-1:0] _tmp_764;
  reg signed [32-1:0] _tmp_765;
  reg signed [32-1:0] _tmp_766;
  reg signed [32-1:0] _tmp_767;
  localparam _tmp_768 = 34;
  wire [_tmp_768-1:0] _tmp_769;
  assign _tmp_769 = _th_comp_size_3 + 32 - 1 >>> 5;
  reg [_tmp_768-1:0] _tmp_770;
  reg [_tmp_768-1:0] _tmp_771;
  reg [_tmp_768-1:0] _tmp_772;
  reg [_tmp_768-1:0] _tmp_773;
  reg [_tmp_768-1:0] _tmp_774;
  reg [_tmp_768-1:0] _tmp_775;
  reg [32-1:0] _mystream_sum_vec18_sink_fsm_82;
  localparam _mystream_sum_vec18_sink_fsm_82_init = 0;
  wire _set_flag_776;
  assign _set_flag_776 = th_comp == 82;
  reg _tmp_777;
  reg _tmp_778;
  reg _tmp_779;
  reg _tmp_780;
  reg _tmp_781;
  reg _tmp_782;
  reg signed [32-1:0] _tmp_783;
  reg signed [32-1:0] _tmp_784;
  reg signed [32-1:0] _tmp_785;
  reg signed [32-1:0] _tmp_786;
  reg signed [32-1:0] _tmp_787;
  reg signed [32-1:0] _tmp_788;
  localparam _tmp_789 = 34;
  wire [_tmp_789-1:0] _tmp_790;
  assign _tmp_790 = _th_comp_size_3 + 32 - 1 >>> 5;
  reg [_tmp_789-1:0] _tmp_791;
  reg [_tmp_789-1:0] _tmp_792;
  reg [_tmp_789-1:0] _tmp_793;
  reg [_tmp_789-1:0] _tmp_794;
  reg [_tmp_789-1:0] _tmp_795;
  reg [_tmp_789-1:0] _tmp_796;
  reg [32-1:0] _mystream_sum_vec19_sink_fsm_83;
  localparam _mystream_sum_vec19_sink_fsm_83_init = 0;
  wire _set_flag_797;
  assign _set_flag_797 = th_comp == 82;
  reg _tmp_798;
  reg _tmp_799;
  reg _tmp_800;
  reg _tmp_801;
  reg _tmp_802;
  reg _tmp_803;
  reg signed [32-1:0] _tmp_804;
  reg signed [32-1:0] _tmp_805;
  reg signed [32-1:0] _tmp_806;
  reg signed [32-1:0] _tmp_807;
  reg signed [32-1:0] _tmp_808;
  reg signed [32-1:0] _tmp_809;
  localparam _tmp_810 = 34;
  wire [_tmp_810-1:0] _tmp_811;
  assign _tmp_811 = _th_comp_size_3 + 32 - 1 >>> 5;
  reg [_tmp_810-1:0] _tmp_812;
  reg [_tmp_810-1:0] _tmp_813;
  reg [_tmp_810-1:0] _tmp_814;
  reg [_tmp_810-1:0] _tmp_815;
  reg [_tmp_810-1:0] _tmp_816;
  reg [_tmp_810-1:0] _tmp_817;
  reg [32-1:0] _mystream_sum_vec20_sink_fsm_84;
  localparam _mystream_sum_vec20_sink_fsm_84_init = 0;
  wire _set_flag_818;
  assign _set_flag_818 = th_comp == 82;
  reg _tmp_819;
  reg _tmp_820;
  reg _tmp_821;
  reg _tmp_822;
  reg _tmp_823;
  reg _tmp_824;
  reg signed [32-1:0] _tmp_825;
  reg signed [32-1:0] _tmp_826;
  reg signed [32-1:0] _tmp_827;
  reg signed [32-1:0] _tmp_828;
  reg signed [32-1:0] _tmp_829;
  reg signed [32-1:0] _tmp_830;
  localparam _tmp_831 = 34;
  wire [_tmp_831-1:0] _tmp_832;
  assign _tmp_832 = _th_comp_size_3 + 32 - 1 >>> 5;
  reg [_tmp_831-1:0] _tmp_833;
  reg [_tmp_831-1:0] _tmp_834;
  reg [_tmp_831-1:0] _tmp_835;
  reg [_tmp_831-1:0] _tmp_836;
  reg [_tmp_831-1:0] _tmp_837;
  reg [_tmp_831-1:0] _tmp_838;
  reg [32-1:0] _mystream_sum_vec21_sink_fsm_85;
  localparam _mystream_sum_vec21_sink_fsm_85_init = 0;
  wire _set_flag_839;
  assign _set_flag_839 = th_comp == 82;
  reg _tmp_840;
  reg _tmp_841;
  reg _tmp_842;
  reg _tmp_843;
  reg _tmp_844;
  reg _tmp_845;
  reg signed [32-1:0] _tmp_846;
  reg signed [32-1:0] _tmp_847;
  reg signed [32-1:0] _tmp_848;
  reg signed [32-1:0] _tmp_849;
  reg signed [32-1:0] _tmp_850;
  reg signed [32-1:0] _tmp_851;
  localparam _tmp_852 = 34;
  wire [_tmp_852-1:0] _tmp_853;
  assign _tmp_853 = _th_comp_size_3 + 32 - 1 >>> 5;
  reg [_tmp_852-1:0] _tmp_854;
  reg [_tmp_852-1:0] _tmp_855;
  reg [_tmp_852-1:0] _tmp_856;
  reg [_tmp_852-1:0] _tmp_857;
  reg [_tmp_852-1:0] _tmp_858;
  reg [_tmp_852-1:0] _tmp_859;
  reg [32-1:0] _mystream_sum_vec22_sink_fsm_86;
  localparam _mystream_sum_vec22_sink_fsm_86_init = 0;
  wire _set_flag_860;
  assign _set_flag_860 = th_comp == 82;
  reg _tmp_861;
  reg _tmp_862;
  reg _tmp_863;
  reg _tmp_864;
  reg _tmp_865;
  reg _tmp_866;
  reg signed [32-1:0] _tmp_867;
  reg signed [32-1:0] _tmp_868;
  reg signed [32-1:0] _tmp_869;
  reg signed [32-1:0] _tmp_870;
  reg signed [32-1:0] _tmp_871;
  reg signed [32-1:0] _tmp_872;
  localparam _tmp_873 = 34;
  wire [_tmp_873-1:0] _tmp_874;
  assign _tmp_874 = _th_comp_size_3 + 32 - 1 >>> 5;
  reg [_tmp_873-1:0] _tmp_875;
  reg [_tmp_873-1:0] _tmp_876;
  reg [_tmp_873-1:0] _tmp_877;
  reg [_tmp_873-1:0] _tmp_878;
  reg [_tmp_873-1:0] _tmp_879;
  reg [_tmp_873-1:0] _tmp_880;
  reg [32-1:0] _mystream_sum_vec23_sink_fsm_87;
  localparam _mystream_sum_vec23_sink_fsm_87_init = 0;
  wire _set_flag_881;
  assign _set_flag_881 = th_comp == 82;
  reg _tmp_882;
  reg _tmp_883;
  reg _tmp_884;
  reg _tmp_885;
  reg _tmp_886;
  reg _tmp_887;
  reg signed [32-1:0] _tmp_888;
  reg signed [32-1:0] _tmp_889;
  reg signed [32-1:0] _tmp_890;
  reg signed [32-1:0] _tmp_891;
  reg signed [32-1:0] _tmp_892;
  reg signed [32-1:0] _tmp_893;
  localparam _tmp_894 = 34;
  wire [_tmp_894-1:0] _tmp_895;
  assign _tmp_895 = _th_comp_size_3 + 32 - 1 >>> 5;
  reg [_tmp_894-1:0] _tmp_896;
  reg [_tmp_894-1:0] _tmp_897;
  reg [_tmp_894-1:0] _tmp_898;
  reg [_tmp_894-1:0] _tmp_899;
  reg [_tmp_894-1:0] _tmp_900;
  reg [_tmp_894-1:0] _tmp_901;
  reg [32-1:0] _mystream_sum_vec24_sink_fsm_88;
  localparam _mystream_sum_vec24_sink_fsm_88_init = 0;
  wire _set_flag_902;
  assign _set_flag_902 = th_comp == 82;
  reg _tmp_903;
  reg _tmp_904;
  reg _tmp_905;
  reg _tmp_906;
  reg _tmp_907;
  reg _tmp_908;
  reg signed [32-1:0] _tmp_909;
  reg signed [32-1:0] _tmp_910;
  reg signed [32-1:0] _tmp_911;
  reg signed [32-1:0] _tmp_912;
  reg signed [32-1:0] _tmp_913;
  reg signed [32-1:0] _tmp_914;
  localparam _tmp_915 = 34;
  wire [_tmp_915-1:0] _tmp_916;
  assign _tmp_916 = _th_comp_size_3 + 32 - 1 >>> 5;
  reg [_tmp_915-1:0] _tmp_917;
  reg [_tmp_915-1:0] _tmp_918;
  reg [_tmp_915-1:0] _tmp_919;
  reg [_tmp_915-1:0] _tmp_920;
  reg [_tmp_915-1:0] _tmp_921;
  reg [_tmp_915-1:0] _tmp_922;
  reg [32-1:0] _mystream_sum_vec25_sink_fsm_89;
  localparam _mystream_sum_vec25_sink_fsm_89_init = 0;
  wire _set_flag_923;
  assign _set_flag_923 = th_comp == 82;
  reg _tmp_924;
  reg _tmp_925;
  reg _tmp_926;
  reg _tmp_927;
  reg _tmp_928;
  reg _tmp_929;
  reg signed [32-1:0] _tmp_930;
  reg signed [32-1:0] _tmp_931;
  reg signed [32-1:0] _tmp_932;
  reg signed [32-1:0] _tmp_933;
  reg signed [32-1:0] _tmp_934;
  reg signed [32-1:0] _tmp_935;
  localparam _tmp_936 = 34;
  wire [_tmp_936-1:0] _tmp_937;
  assign _tmp_937 = _th_comp_size_3 + 32 - 1 >>> 5;
  reg [_tmp_936-1:0] _tmp_938;
  reg [_tmp_936-1:0] _tmp_939;
  reg [_tmp_936-1:0] _tmp_940;
  reg [_tmp_936-1:0] _tmp_941;
  reg [_tmp_936-1:0] _tmp_942;
  reg [_tmp_936-1:0] _tmp_943;
  reg [32-1:0] _mystream_sum_vec26_sink_fsm_90;
  localparam _mystream_sum_vec26_sink_fsm_90_init = 0;
  wire _set_flag_944;
  assign _set_flag_944 = th_comp == 82;
  reg _tmp_945;
  reg _tmp_946;
  reg _tmp_947;
  reg _tmp_948;
  reg _tmp_949;
  reg _tmp_950;
  reg signed [32-1:0] _tmp_951;
  reg signed [32-1:0] _tmp_952;
  reg signed [32-1:0] _tmp_953;
  reg signed [32-1:0] _tmp_954;
  reg signed [32-1:0] _tmp_955;
  reg signed [32-1:0] _tmp_956;
  localparam _tmp_957 = 34;
  wire [_tmp_957-1:0] _tmp_958;
  assign _tmp_958 = _th_comp_size_3 + 32 - 1 >>> 5;
  reg [_tmp_957-1:0] _tmp_959;
  reg [_tmp_957-1:0] _tmp_960;
  reg [_tmp_957-1:0] _tmp_961;
  reg [_tmp_957-1:0] _tmp_962;
  reg [_tmp_957-1:0] _tmp_963;
  reg [_tmp_957-1:0] _tmp_964;
  reg [32-1:0] _mystream_sum_vec27_sink_fsm_91;
  localparam _mystream_sum_vec27_sink_fsm_91_init = 0;
  wire _set_flag_965;
  assign _set_flag_965 = th_comp == 82;
  reg _tmp_966;
  reg _tmp_967;
  reg _tmp_968;
  reg _tmp_969;
  reg _tmp_970;
  reg _tmp_971;
  reg signed [32-1:0] _tmp_972;
  reg signed [32-1:0] _tmp_973;
  reg signed [32-1:0] _tmp_974;
  reg signed [32-1:0] _tmp_975;
  reg signed [32-1:0] _tmp_976;
  reg signed [32-1:0] _tmp_977;
  localparam _tmp_978 = 34;
  wire [_tmp_978-1:0] _tmp_979;
  assign _tmp_979 = _th_comp_size_3 + 32 - 1 >>> 5;
  reg [_tmp_978-1:0] _tmp_980;
  reg [_tmp_978-1:0] _tmp_981;
  reg [_tmp_978-1:0] _tmp_982;
  reg [_tmp_978-1:0] _tmp_983;
  reg [_tmp_978-1:0] _tmp_984;
  reg [_tmp_978-1:0] _tmp_985;
  reg [32-1:0] _mystream_sum_vec28_sink_fsm_92;
  localparam _mystream_sum_vec28_sink_fsm_92_init = 0;
  wire _set_flag_986;
  assign _set_flag_986 = th_comp == 82;
  reg _tmp_987;
  reg _tmp_988;
  reg _tmp_989;
  reg _tmp_990;
  reg _tmp_991;
  reg _tmp_992;
  reg signed [32-1:0] _tmp_993;
  reg signed [32-1:0] _tmp_994;
  reg signed [32-1:0] _tmp_995;
  reg signed [32-1:0] _tmp_996;
  reg signed [32-1:0] _tmp_997;
  reg signed [32-1:0] _tmp_998;
  localparam _tmp_999 = 34;
  wire [_tmp_999-1:0] _tmp_1000;
  assign _tmp_1000 = _th_comp_size_3 + 32 - 1 >>> 5;
  reg [_tmp_999-1:0] _tmp_1001;
  reg [_tmp_999-1:0] _tmp_1002;
  reg [_tmp_999-1:0] _tmp_1003;
  reg [_tmp_999-1:0] _tmp_1004;
  reg [_tmp_999-1:0] _tmp_1005;
  reg [_tmp_999-1:0] _tmp_1006;
  reg [32-1:0] _mystream_sum_vec29_sink_fsm_93;
  localparam _mystream_sum_vec29_sink_fsm_93_init = 0;
  wire _set_flag_1007;
  assign _set_flag_1007 = th_comp == 82;
  reg _tmp_1008;
  reg _tmp_1009;
  reg _tmp_1010;
  reg _tmp_1011;
  reg _tmp_1012;
  reg _tmp_1013;
  reg signed [32-1:0] _tmp_1014;
  reg signed [32-1:0] _tmp_1015;
  reg signed [32-1:0] _tmp_1016;
  reg signed [32-1:0] _tmp_1017;
  reg signed [32-1:0] _tmp_1018;
  reg signed [32-1:0] _tmp_1019;
  localparam _tmp_1020 = 34;
  wire [_tmp_1020-1:0] _tmp_1021;
  assign _tmp_1021 = _th_comp_size_3 + 32 - 1 >>> 5;
  reg [_tmp_1020-1:0] _tmp_1022;
  reg [_tmp_1020-1:0] _tmp_1023;
  reg [_tmp_1020-1:0] _tmp_1024;
  reg [_tmp_1020-1:0] _tmp_1025;
  reg [_tmp_1020-1:0] _tmp_1026;
  reg [_tmp_1020-1:0] _tmp_1027;
  reg [32-1:0] _mystream_sum_vec30_sink_fsm_94;
  localparam _mystream_sum_vec30_sink_fsm_94_init = 0;
  wire _set_flag_1028;
  assign _set_flag_1028 = th_comp == 82;
  reg _tmp_1029;
  reg _tmp_1030;
  reg _tmp_1031;
  reg _tmp_1032;
  reg _tmp_1033;
  reg _tmp_1034;
  reg signed [32-1:0] _tmp_1035;
  reg signed [32-1:0] _tmp_1036;
  reg signed [32-1:0] _tmp_1037;
  reg signed [32-1:0] _tmp_1038;
  reg signed [32-1:0] _tmp_1039;
  reg signed [32-1:0] _tmp_1040;
  localparam _tmp_1041 = 34;
  wire [_tmp_1041-1:0] _tmp_1042;
  assign _tmp_1042 = _th_comp_size_3 + 32 - 1 >>> 5;
  reg [_tmp_1041-1:0] _tmp_1043;
  reg [_tmp_1041-1:0] _tmp_1044;
  reg [_tmp_1041-1:0] _tmp_1045;
  reg [_tmp_1041-1:0] _tmp_1046;
  reg [_tmp_1041-1:0] _tmp_1047;
  reg [_tmp_1041-1:0] _tmp_1048;
  reg [32-1:0] _mystream_sum_vec31_sink_fsm_95;
  localparam _mystream_sum_vec31_sink_fsm_95_init = 0;
  wire _set_flag_1049;
  assign _set_flag_1049 = th_comp == 84;
  assign _mystream_run_flag = (_set_flag_1049)? 1 : 0;
  reg _tmp_1050;
  reg _tmp_1051;
  reg _tmp_1052;
  reg _tmp_1053;
  reg _tmp_1054;
  reg _tmp_1055;
  reg [1-1:0] __variable_wdata_130;
  assign mystream__reduce_reset_data = __variable_wdata_130;
  reg _tmp_1056;
  reg _tmp_1057;
  reg _tmp_1058;
  reg _tmp_1059;
  assign _mystream_source_stop = _mystream_stream_oready && (_mystream_a0_idle && _mystream_a1_idle && _mystream_a10_idle && _mystream_a11_idle && _mystream_a12_idle && _mystream_a13_idle && _mystream_a14_idle && _mystream_a15_idle && _mystream_a16_idle && _mystream_a17_idle && _mystream_a18_idle && _mystream_a19_idle && _mystream_a2_idle && _mystream_a20_idle && _mystream_a21_idle && _mystream_a22_idle && _mystream_a23_idle && _mystream_a24_idle && _mystream_a25_idle && _mystream_a26_idle && _mystream_a27_idle && _mystream_a28_idle && _mystream_a29_idle && _mystream_a3_idle && _mystream_a30_idle && _mystream_a31_idle && _mystream_a4_idle && _mystream_a5_idle && _mystream_a6_idle && _mystream_a7_idle && _mystream_a8_idle && _mystream_a9_idle && _mystream_b0_idle && _mystream_b1_idle && _mystream_b10_idle && _mystream_b11_idle && _mystream_b12_idle && _mystream_b13_idle && _mystream_b14_idle && _mystream_b15_idle && _mystream_b16_idle && _mystream_b17_idle && _mystream_b18_idle && _mystream_b19_idle && _mystream_b2_idle && _mystream_b20_idle && _mystream_b21_idle && _mystream_b22_idle && _mystream_b23_idle && _mystream_b24_idle && _mystream_b25_idle && _mystream_b26_idle && _mystream_b27_idle && _mystream_b28_idle && _mystream_b29_idle && _mystream_b3_idle && _mystream_b30_idle && _mystream_b31_idle && _mystream_b4_idle && _mystream_b5_idle && _mystream_b6_idle && _mystream_b7_idle && _mystream_b8_idle && _mystream_b9_idle && _mystream_bias0_idle && _mystream_bias1_idle && _mystream_bias10_idle && _mystream_bias11_idle && _mystream_bias12_idle && _mystream_bias13_idle && _mystream_bias14_idle && _mystream_bias15_idle && _mystream_bias16_idle && _mystream_bias17_idle && _mystream_bias18_idle && _mystream_bias19_idle && _mystream_bias2_idle && _mystream_bias20_idle && _mystream_bias21_idle && _mystream_bias22_idle && _mystream_bias23_idle && _mystream_bias24_idle && _mystream_bias25_idle && _mystream_bias26_idle && _mystream_bias27_idle && _mystream_bias28_idle && _mystream_bias29_idle && _mystream_bias3_idle && _mystream_bias30_idle && _mystream_bias31_idle && _mystream_bias4_idle && _mystream_bias5_idle && _mystream_bias6_idle && _mystream_bias7_idle && _mystream_bias8_idle && _mystream_bias9_idle && (_mystream_fsm == 3));
  localparam _tmp_1060 = 1;
  wire [_tmp_1060-1:0] _tmp_1061;
  assign _tmp_1061 = _mystream_a0_idle && _mystream_a1_idle && _mystream_a10_idle && _mystream_a11_idle && _mystream_a12_idle && _mystream_a13_idle && _mystream_a14_idle && _mystream_a15_idle && _mystream_a16_idle && _mystream_a17_idle && _mystream_a18_idle && _mystream_a19_idle && _mystream_a2_idle && _mystream_a20_idle && _mystream_a21_idle && _mystream_a22_idle && _mystream_a23_idle && _mystream_a24_idle && _mystream_a25_idle && _mystream_a26_idle && _mystream_a27_idle && _mystream_a28_idle && _mystream_a29_idle && _mystream_a3_idle && _mystream_a30_idle && _mystream_a31_idle && _mystream_a4_idle && _mystream_a5_idle && _mystream_a6_idle && _mystream_a7_idle && _mystream_a8_idle && _mystream_a9_idle && _mystream_b0_idle && _mystream_b1_idle && _mystream_b10_idle && _mystream_b11_idle && _mystream_b12_idle && _mystream_b13_idle && _mystream_b14_idle && _mystream_b15_idle && _mystream_b16_idle && _mystream_b17_idle && _mystream_b18_idle && _mystream_b19_idle && _mystream_b2_idle && _mystream_b20_idle && _mystream_b21_idle && _mystream_b22_idle && _mystream_b23_idle && _mystream_b24_idle && _mystream_b25_idle && _mystream_b26_idle && _mystream_b27_idle && _mystream_b28_idle && _mystream_b29_idle && _mystream_b3_idle && _mystream_b30_idle && _mystream_b31_idle && _mystream_b4_idle && _mystream_b5_idle && _mystream_b6_idle && _mystream_b7_idle && _mystream_b8_idle && _mystream_b9_idle && _mystream_bias0_idle && _mystream_bias1_idle && _mystream_bias10_idle && _mystream_bias11_idle && _mystream_bias12_idle && _mystream_bias13_idle && _mystream_bias14_idle && _mystream_bias15_idle && _mystream_bias16_idle && _mystream_bias17_idle && _mystream_bias18_idle && _mystream_bias19_idle && _mystream_bias2_idle && _mystream_bias20_idle && _mystream_bias21_idle && _mystream_bias22_idle && _mystream_bias23_idle && _mystream_bias24_idle && _mystream_bias25_idle && _mystream_bias26_idle && _mystream_bias27_idle && _mystream_bias28_idle && _mystream_bias29_idle && _mystream_bias3_idle && _mystream_bias30_idle && _mystream_bias31_idle && _mystream_bias4_idle && _mystream_bias5_idle && _mystream_bias6_idle && _mystream_bias7_idle && _mystream_bias8_idle && _mystream_bias9_idle && (_mystream_fsm == 3);
  reg [_tmp_1060-1:0] _tmp_1062;
  localparam _tmp_1063 = 1;
  wire [_tmp_1063-1:0] _tmp_1064;
  assign _tmp_1064 = _mystream_a0_idle && _mystream_a1_idle && _mystream_a10_idle && _mystream_a11_idle && _mystream_a12_idle && _mystream_a13_idle && _mystream_a14_idle && _mystream_a15_idle && _mystream_a16_idle && _mystream_a17_idle && _mystream_a18_idle && _mystream_a19_idle && _mystream_a2_idle && _mystream_a20_idle && _mystream_a21_idle && _mystream_a22_idle && _mystream_a23_idle && _mystream_a24_idle && _mystream_a25_idle && _mystream_a26_idle && _mystream_a27_idle && _mystream_a28_idle && _mystream_a29_idle && _mystream_a3_idle && _mystream_a30_idle && _mystream_a31_idle && _mystream_a4_idle && _mystream_a5_idle && _mystream_a6_idle && _mystream_a7_idle && _mystream_a8_idle && _mystream_a9_idle && _mystream_b0_idle && _mystream_b1_idle && _mystream_b10_idle && _mystream_b11_idle && _mystream_b12_idle && _mystream_b13_idle && _mystream_b14_idle && _mystream_b15_idle && _mystream_b16_idle && _mystream_b17_idle && _mystream_b18_idle && _mystream_b19_idle && _mystream_b2_idle && _mystream_b20_idle && _mystream_b21_idle && _mystream_b22_idle && _mystream_b23_idle && _mystream_b24_idle && _mystream_b25_idle && _mystream_b26_idle && _mystream_b27_idle && _mystream_b28_idle && _mystream_b29_idle && _mystream_b3_idle && _mystream_b30_idle && _mystream_b31_idle && _mystream_b4_idle && _mystream_b5_idle && _mystream_b6_idle && _mystream_b7_idle && _mystream_b8_idle && _mystream_b9_idle && _mystream_bias0_idle && _mystream_bias1_idle && _mystream_bias10_idle && _mystream_bias11_idle && _mystream_bias12_idle && _mystream_bias13_idle && _mystream_bias14_idle && _mystream_bias15_idle && _mystream_bias16_idle && _mystream_bias17_idle && _mystream_bias18_idle && _mystream_bias19_idle && _mystream_bias2_idle && _mystream_bias20_idle && _mystream_bias21_idle && _mystream_bias22_idle && _mystream_bias23_idle && _mystream_bias24_idle && _mystream_bias25_idle && _mystream_bias26_idle && _mystream_bias27_idle && _mystream_bias28_idle && _mystream_bias29_idle && _mystream_bias3_idle && _mystream_bias30_idle && _mystream_bias31_idle && _mystream_bias4_idle && _mystream_bias5_idle && _mystream_bias6_idle && _mystream_bias7_idle && _mystream_bias8_idle && _mystream_bias9_idle && (_mystream_fsm == 3);
  reg [_tmp_1063-1:0] _tmp_1065;
  reg _tmp_1066;
  reg _tmp_1067;
  reg _tmp_1068;
  reg _tmp_1069;
  reg _tmp_1070;
  reg _tmp_1071;
  assign _mystream_sink_start = _tmp_1071;
  reg _tmp_1072;
  reg _tmp_1073;
  reg _tmp_1074;
  reg _tmp_1075;
  reg _tmp_1076;
  reg _tmp_1077;
  assign _mystream_sink_stop = _tmp_1077;
  reg _tmp_1078;
  reg _tmp_1079;
  reg _tmp_1080;
  reg _tmp_1081;
  reg _tmp_1082;
  reg _tmp_1083;
  assign _mystream_sink_busy = _tmp_1083;
  reg _tmp_1084;
  assign _mystream_busy = _mystream_source_busy || _mystream_sink_busy || _mystream_busy_reg;
  reg signed [32-1:0] _th_comp_exec_time_7;
  wire [32-1:0] mask_addr_shifted_1085;
  assign mask_addr_shifted_1085 = 0 + (_th_comp_size_0 << 2) >> 2;
  wire [32-1:0] mask_addr_masked_1086;
  assign mask_addr_masked_1086 = mask_addr_shifted_1085 << 2;
  reg [32-1:0] _myaxi_read_data_fsm;
  localparam _myaxi_read_data_fsm_init = 0;
  reg [32-1:0] write_burst_fsm_2;
  localparam write_burst_fsm_2_init = 0;
  reg [20-1:0] write_burst_addr_1087;
  reg [20-1:0] write_burst_stride_1088;
  reg [33-1:0] write_burst_length_1089;
  reg write_burst_done_1090;
  assign ram_x_0_wdata = ((write_burst_fsm_2 == 1) && myaxi_rvalid)? myaxi_rdata : 'hx;
  assign ram_x_0_wenable = ((write_burst_fsm_2 == 1) && myaxi_rvalid)? 1'd1 : 0;
  wire [32-1:0] mask_addr_shifted_1091;
  assign mask_addr_shifted_1091 = _th_comp_offset_b_1 + (_th_comp_size_0 << 2) >> 2;
  wire [32-1:0] mask_addr_masked_1092;
  assign mask_addr_masked_1092 = mask_addr_shifted_1091 << 2;
  reg [32-1:0] write_burst_fsm_3;
  localparam write_burst_fsm_3_init = 0;
  reg [20-1:0] write_burst_addr_1093;
  reg [20-1:0] write_burst_stride_1094;
  reg [33-1:0] write_burst_length_1095;
  reg write_burst_done_1096;
  assign ram_y_0_wdata = ((write_burst_fsm_3 == 1) && myaxi_rvalid)? myaxi_rdata : 'hx;
  assign ram_y_0_wenable = ((write_burst_fsm_3 == 1) && myaxi_rvalid)? 1'd1 : 0;
  reg signed [32-1:0] _th_comp_size_8;
  reg signed [32-1:0] _th_comp_offset_9;
  reg signed [32-1:0] _th_comp_sum_10;
  reg signed [32-1:0] _th_comp_i_11;
  assign ram_x_0_addr = (th_comp == 99)? _th_comp_i_11 + _th_comp_offset_9 : 
                        ((write_burst_fsm_2 == 1) && myaxi_rvalid)? write_burst_addr_1087 : 'hx;
  assign ram_x_0_enable = (th_comp == 99)? 1'd1 : 
                          ((write_burst_fsm_2 == 1) && myaxi_rvalid)? 1'd1 : 0;
  localparam _tmp_1097 = 1;
  wire [_tmp_1097-1:0] _tmp_1098;
  assign _tmp_1098 = th_comp == 99;
  reg [_tmp_1097-1:0] __tmp_1098_1;
  reg signed [32-1:0] read_rdata_1099;
  reg signed [32-1:0] _th_comp_a_12;
  assign ram_y_0_addr = (th_comp == 101)? _th_comp_i_11 + _th_comp_offset_9 : 
                        ((write_burst_fsm_3 == 1) && myaxi_rvalid)? write_burst_addr_1093 : 'hx;
  assign ram_y_0_enable = (th_comp == 101)? 1'd1 : 
                          ((write_burst_fsm_3 == 1) && myaxi_rvalid)? 1'd1 : 0;
  localparam _tmp_1100 = 1;
  wire [_tmp_1100-1:0] _tmp_1101;
  assign _tmp_1101 = th_comp == 101;
  reg [_tmp_1100-1:0] __tmp_1101_1;
  reg signed [32-1:0] read_rdata_1102;
  reg signed [32-1:0] _th_comp_b_13;
  assign ram_z_0_wdata = (th_comp == 104)? _th_comp_sum_10 : 'hx;
  assign ram_z_0_wenable = (th_comp == 104)? 1'd1 : 0;
  wire [32-1:0] mask_addr_shifted_1103;
  assign mask_addr_shifted_1103 = 2048 >> 2;
  wire [32-1:0] mask_addr_masked_1104;
  assign mask_addr_masked_1104 = mask_addr_shifted_1103 << 2;
  reg [32-1:0] _myaxi_write_req_fsm;
  localparam _myaxi_write_req_fsm_init = 0;
  reg [33-1:0] _myaxi_write_cur_global_size;
  reg _myaxi_write_cont;
  wire [8-1:0] pack_write_req_op_sel_1105;
  wire [32-1:0] pack_write_req_local_addr_1106;
  wire [32-1:0] pack_write_req_local_stride_1107;
  wire [33-1:0] pack_write_req_size_1108;
  wire [32-1:0] pack_write_req_local_blocksize_1109;
  assign pack_write_req_op_sel_1105 = _myaxi_write_op_sel;
  assign pack_write_req_local_addr_1106 = _myaxi_write_local_addr;
  assign pack_write_req_local_stride_1107 = _myaxi_write_local_stride;
  assign pack_write_req_size_1108 = _myaxi_write_local_size;
  assign pack_write_req_local_blocksize_1109 = _myaxi_write_local_blocksize;
  wire [137-1:0] pack_write_req_packed_1110;
  assign pack_write_req_packed_1110 = { pack_write_req_op_sel_1105, pack_write_req_local_addr_1106, pack_write_req_local_stride_1107, pack_write_req_size_1108, pack_write_req_local_blocksize_1109 };
  localparam _tmp_1111 = 1;
  wire [_tmp_1111-1:0] _tmp_1112;
  assign _tmp_1112 = !_myaxi_write_req_fifo_almost_full;
  reg [_tmp_1111-1:0] __tmp_1112_1;
  wire [32-1:0] mask_addr_shifted_1113;
  assign mask_addr_shifted_1113 = _myaxi_write_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_1114;
  assign mask_addr_masked_1114 = mask_addr_shifted_1113 << 2;
  wire [32-1:0] mask_addr_shifted_1115;
  assign mask_addr_shifted_1115 = _myaxi_write_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_1116;
  assign mask_addr_masked_1116 = mask_addr_shifted_1115 << 2;
  wire [32-1:0] mask_addr_shifted_1117;
  assign mask_addr_shifted_1117 = _myaxi_write_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_1118;
  assign mask_addr_masked_1118 = mask_addr_shifted_1117 << 2;
  wire [32-1:0] mask_addr_shifted_1119;
  assign mask_addr_shifted_1119 = _myaxi_write_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_1120;
  assign mask_addr_masked_1120 = mask_addr_shifted_1119 << 2;
  wire [32-1:0] mask_addr_shifted_1121;
  assign mask_addr_shifted_1121 = _myaxi_write_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_1122;
  assign mask_addr_masked_1122 = mask_addr_shifted_1121 << 2;
  wire [32-1:0] mask_addr_shifted_1123;
  assign mask_addr_shifted_1123 = _myaxi_write_global_addr >> 2;
  wire [32-1:0] mask_addr_masked_1124;
  assign mask_addr_masked_1124 = mask_addr_shifted_1123 << 2;
  wire [8-1:0] pack_write_req_op_sel_1125;
  wire [32-1:0] pack_write_req_local_addr_1126;
  wire [32-1:0] pack_write_req_local_stride_1127;
  wire [33-1:0] pack_write_req_size_1128;
  wire [32-1:0] pack_write_req_local_blocksize_1129;
  assign pack_write_req_op_sel_1125 = _myaxi_write_op_sel;
  assign pack_write_req_local_addr_1126 = _myaxi_write_local_addr;
  assign pack_write_req_local_stride_1127 = _myaxi_write_local_stride;
  assign pack_write_req_size_1128 = _myaxi_write_cur_global_size;
  assign pack_write_req_local_blocksize_1129 = _myaxi_write_local_blocksize;
  wire [137-1:0] pack_write_req_packed_1130;
  assign pack_write_req_packed_1130 = { pack_write_req_op_sel_1125, pack_write_req_local_addr_1126, pack_write_req_local_stride_1127, pack_write_req_size_1128, pack_write_req_local_blocksize_1129 };
  assign _myaxi_write_req_fifo_wdata = ((_myaxi_write_req_fsm == 1) && !_myaxi_write_req_fifo_almost_full && (myaxi_awready || !myaxi_awvalid) && (outstanding_wcount_0 < 6))? pack_write_req_packed_1130 : 
                                       ((_myaxi_write_req_fsm == 0) && _myaxi_write_start && !_myaxi_write_req_fifo_almost_full)? pack_write_req_packed_1110 : 'hx;
  assign _myaxi_write_req_fifo_enq = ((_myaxi_write_req_fsm == 1) && !_myaxi_write_req_fifo_almost_full && (myaxi_awready || !myaxi_awvalid) && (outstanding_wcount_0 < 6))? (_myaxi_write_req_fsm == 1) && !_myaxi_write_req_fifo_almost_full && (myaxi_awready || !myaxi_awvalid) && (outstanding_wcount_0 < 6) && !_myaxi_write_req_fifo_almost_full : 
                                     ((_myaxi_write_req_fsm == 0) && _myaxi_write_start && !_myaxi_write_req_fifo_almost_full)? (_myaxi_write_req_fsm == 0) && _myaxi_write_start && !_myaxi_write_req_fifo_almost_full && !_myaxi_write_req_fifo_almost_full : 0;
  localparam _tmp_1131 = 1;
  wire [_tmp_1131-1:0] _tmp_1132;
  assign _tmp_1132 = !_myaxi_write_req_fifo_almost_full;
  reg [_tmp_1131-1:0] __tmp_1132_1;
  reg _myaxi_cond_1_1;
  reg [32-1:0] _myaxi_write_data_fsm;
  localparam _myaxi_write_data_fsm_init = 0;
  reg [32-1:0] read_burst_fsm_4;
  localparam read_burst_fsm_4_init = 0;
  reg [20-1:0] read_burst_addr_1133;
  reg [20-1:0] read_burst_stride_1134;
  reg [33-1:0] read_burst_length_1135;
  reg read_burst_rvalid_1136;
  reg read_burst_rlast_1137;
  assign ram_z_0_addr = ((read_burst_fsm_4 == 1) && (!read_burst_rvalid_1136 || (myaxi_wready || !myaxi_wvalid) && (_myaxi_write_size_buf > 0)))? read_burst_addr_1133 : 
                        (th_comp == 104)? _th_comp_i_11 + _th_comp_offset_9 : 'hx;
  assign ram_z_0_enable = ((read_burst_fsm_4 == 1) && (!read_burst_rvalid_1136 || (myaxi_wready || !myaxi_wvalid) && (_myaxi_write_size_buf > 0)))? 1'd1 : 
                          (th_comp == 104)? 1'd1 : 0;
  localparam _tmp_1138 = 1;
  wire [_tmp_1138-1:0] _tmp_1139;
  assign _tmp_1139 = (read_burst_fsm_4 == 1) && (!read_burst_rvalid_1136 || (myaxi_wready || !myaxi_wvalid) && (_myaxi_write_size_buf > 0));
  reg [_tmp_1138-1:0] __tmp_1139_1;
  wire [32-1:0] read_burst_rdata_1140;
  assign read_burst_rdata_1140 = ram_z_0_rdata;
  assign _myaxi_write_req_fifo_deq = ((_myaxi_write_data_fsm == 2) && (!_myaxi_write_req_fifo_empty && (_myaxi_write_size_buf == 0)) && !_myaxi_write_req_fifo_empty)? 1 : 
                                     ((_myaxi_write_data_fsm == 0) && (_myaxi_write_data_idle && !_myaxi_write_req_fifo_empty && (_myaxi_write_op_sel_fifo == 1)) && !_myaxi_write_req_fifo_empty)? 1 : 0;
  reg _myaxi_cond_2_1;
  wire [32-1:0] _dma_read_packed_high_local_size_1141;
  assign _dma_read_packed_high_local_size_1141 = _th_comp_size_0 >> 5;
  wire [5-1:0] _dma_read_packed_low_local_size_1142;
  assign _dma_read_packed_low_local_size_1142 = _th_comp_size_0 & { 5{ 1'd1 } };
  wire [32-1:0] _dma_read_packed_local_packed_size_1143;
  assign _dma_read_packed_local_packed_size_1143 = (_dma_read_packed_low_local_size_1142 > 0)? _dma_read_packed_high_local_size_1141 + 1 : _dma_read_packed_high_local_size_1141;
  wire [32-1:0] mask_addr_shifted_1144;
  assign mask_addr_shifted_1144 = 2048 >> 2;
  wire [32-1:0] mask_addr_masked_1145;
  assign mask_addr_masked_1145 = mask_addr_shifted_1144 << 2;
  assign _myaxi_read_req_fifo_deq = ((_myaxi_read_data_narrow_fsm == 0) && (_myaxi_read_data_idle && !_myaxi_read_req_fifo_empty && (_myaxi_read_op_sel_fifo == 5)) && !_myaxi_read_req_fifo_empty)? 1 : 
                                    ((_myaxi_read_data_fsm == 0) && (_myaxi_read_data_idle && !_myaxi_read_req_fifo_empty && (_myaxi_read_op_sel_fifo == 4)) && !_myaxi_read_req_fifo_empty)? 1 : 
                                    ((_myaxi_read_data_fsm == 0) && (_myaxi_read_data_idle && !_myaxi_read_req_fifo_empty && (_myaxi_read_op_sel_fifo == 3)) && !_myaxi_read_req_fifo_empty)? 1 : 
                                    ((_myaxi_read_data_narrow_fsm == 0) && (_myaxi_read_data_idle && !_myaxi_read_req_fifo_empty && (_myaxi_read_op_sel_fifo == 2)) && !_myaxi_read_req_fifo_empty)? 1 : 
                                    ((_myaxi_read_data_narrow_fsm == 0) && (_myaxi_read_data_idle && !_myaxi_read_req_fifo_empty && (_myaxi_read_op_sel_fifo == 1)) && !_myaxi_read_req_fifo_empty)? 1 : 0;
  reg [1024-1:0] _myaxi_read_narrow_wdata_1146;
  reg _myaxi_read_narrow_wvalid_1147;
  reg [5-1:0] _myaxi_read_narrow_count_1148;
  reg [32-1:0] write_burst_packed_fsm_5;
  localparam write_burst_packed_fsm_5_init = 0;
  reg [25-1:0] write_burst_packed_addr_1149;
  reg [25-1:0] write_burst_packed_stride_1150;
  reg [33-1:0] write_burst_packed_length_1151;
  reg write_burst_packed_done_1152;
  wire [20-1:0] write_burst_packed_ram_addr_1153;
  assign write_burst_packed_ram_addr_1153 = write_burst_packed_addr_1149 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_1154;
  assign write_burst_packed_ram_wdata_1154 = _myaxi_read_narrow_wdata_1146 >> 0;
  assign ram_c_0_0_wdata = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_wdata_1154 : 
                           (_mystream_stream_oready && _mystream_sum_vec0_sink_wenable && (_mystream_sum_vec0_sink_sel == 65))? _mystream_sum_vec0_sink_wdata : 'hx;
  assign ram_c_0_0_wenable = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                             (_mystream_stream_oready && _mystream_sum_vec0_sink_wenable && (_mystream_sum_vec0_sink_sel == 65))? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_1155;
  assign write_burst_packed_ram_addr_1155 = write_burst_packed_addr_1149 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_1156;
  assign write_burst_packed_ram_wdata_1156 = _myaxi_read_narrow_wdata_1146 >> 32;
  assign ram_c_1_0_wdata = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_wdata_1156 : 
                           (_mystream_stream_oready && _mystream_sum_vec1_sink_wenable && (_mystream_sum_vec1_sink_sel == 66))? _mystream_sum_vec1_sink_wdata : 'hx;
  assign ram_c_1_0_wenable = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                             (_mystream_stream_oready && _mystream_sum_vec1_sink_wenable && (_mystream_sum_vec1_sink_sel == 66))? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_1157;
  assign write_burst_packed_ram_addr_1157 = write_burst_packed_addr_1149 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_1158;
  assign write_burst_packed_ram_wdata_1158 = _myaxi_read_narrow_wdata_1146 >> 64;
  assign ram_c_2_0_wdata = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_wdata_1158 : 
                           (_mystream_stream_oready && _mystream_sum_vec2_sink_wenable && (_mystream_sum_vec2_sink_sel == 67))? _mystream_sum_vec2_sink_wdata : 'hx;
  assign ram_c_2_0_wenable = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                             (_mystream_stream_oready && _mystream_sum_vec2_sink_wenable && (_mystream_sum_vec2_sink_sel == 67))? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_1159;
  assign write_burst_packed_ram_addr_1159 = write_burst_packed_addr_1149 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_1160;
  assign write_burst_packed_ram_wdata_1160 = _myaxi_read_narrow_wdata_1146 >> 96;
  assign ram_c_3_0_wdata = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_wdata_1160 : 
                           (_mystream_stream_oready && _mystream_sum_vec3_sink_wenable && (_mystream_sum_vec3_sink_sel == 68))? _mystream_sum_vec3_sink_wdata : 'hx;
  assign ram_c_3_0_wenable = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                             (_mystream_stream_oready && _mystream_sum_vec3_sink_wenable && (_mystream_sum_vec3_sink_sel == 68))? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_1161;
  assign write_burst_packed_ram_addr_1161 = write_burst_packed_addr_1149 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_1162;
  assign write_burst_packed_ram_wdata_1162 = _myaxi_read_narrow_wdata_1146 >> 128;
  assign ram_c_4_0_wdata = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_wdata_1162 : 
                           (_mystream_stream_oready && _mystream_sum_vec4_sink_wenable && (_mystream_sum_vec4_sink_sel == 69))? _mystream_sum_vec4_sink_wdata : 'hx;
  assign ram_c_4_0_wenable = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                             (_mystream_stream_oready && _mystream_sum_vec4_sink_wenable && (_mystream_sum_vec4_sink_sel == 69))? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_1163;
  assign write_burst_packed_ram_addr_1163 = write_burst_packed_addr_1149 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_1164;
  assign write_burst_packed_ram_wdata_1164 = _myaxi_read_narrow_wdata_1146 >> 160;
  assign ram_c_5_0_wdata = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_wdata_1164 : 
                           (_mystream_stream_oready && _mystream_sum_vec5_sink_wenable && (_mystream_sum_vec5_sink_sel == 70))? _mystream_sum_vec5_sink_wdata : 'hx;
  assign ram_c_5_0_wenable = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                             (_mystream_stream_oready && _mystream_sum_vec5_sink_wenable && (_mystream_sum_vec5_sink_sel == 70))? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_1165;
  assign write_burst_packed_ram_addr_1165 = write_burst_packed_addr_1149 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_1166;
  assign write_burst_packed_ram_wdata_1166 = _myaxi_read_narrow_wdata_1146 >> 192;
  assign ram_c_6_0_wdata = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_wdata_1166 : 
                           (_mystream_stream_oready && _mystream_sum_vec6_sink_wenable && (_mystream_sum_vec6_sink_sel == 71))? _mystream_sum_vec6_sink_wdata : 'hx;
  assign ram_c_6_0_wenable = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                             (_mystream_stream_oready && _mystream_sum_vec6_sink_wenable && (_mystream_sum_vec6_sink_sel == 71))? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_1167;
  assign write_burst_packed_ram_addr_1167 = write_burst_packed_addr_1149 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_1168;
  assign write_burst_packed_ram_wdata_1168 = _myaxi_read_narrow_wdata_1146 >> 224;
  assign ram_c_7_0_wdata = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_wdata_1168 : 
                           (_mystream_stream_oready && _mystream_sum_vec7_sink_wenable && (_mystream_sum_vec7_sink_sel == 72))? _mystream_sum_vec7_sink_wdata : 'hx;
  assign ram_c_7_0_wenable = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                             (_mystream_stream_oready && _mystream_sum_vec7_sink_wenable && (_mystream_sum_vec7_sink_sel == 72))? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_1169;
  assign write_burst_packed_ram_addr_1169 = write_burst_packed_addr_1149 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_1170;
  assign write_burst_packed_ram_wdata_1170 = _myaxi_read_narrow_wdata_1146 >> 256;
  assign ram_c_8_0_wdata = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_wdata_1170 : 
                           (_mystream_stream_oready && _mystream_sum_vec8_sink_wenable && (_mystream_sum_vec8_sink_sel == 73))? _mystream_sum_vec8_sink_wdata : 'hx;
  assign ram_c_8_0_wenable = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                             (_mystream_stream_oready && _mystream_sum_vec8_sink_wenable && (_mystream_sum_vec8_sink_sel == 73))? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_1171;
  assign write_burst_packed_ram_addr_1171 = write_burst_packed_addr_1149 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_1172;
  assign write_burst_packed_ram_wdata_1172 = _myaxi_read_narrow_wdata_1146 >> 288;
  assign ram_c_9_0_wdata = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_wdata_1172 : 
                           (_mystream_stream_oready && _mystream_sum_vec9_sink_wenable && (_mystream_sum_vec9_sink_sel == 74))? _mystream_sum_vec9_sink_wdata : 'hx;
  assign ram_c_9_0_wenable = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                             (_mystream_stream_oready && _mystream_sum_vec9_sink_wenable && (_mystream_sum_vec9_sink_sel == 74))? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_1173;
  assign write_burst_packed_ram_addr_1173 = write_burst_packed_addr_1149 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_1174;
  assign write_burst_packed_ram_wdata_1174 = _myaxi_read_narrow_wdata_1146 >> 320;
  assign ram_c_10_0_wdata = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_wdata_1174 : 
                            (_mystream_stream_oready && _mystream_sum_vec10_sink_wenable && (_mystream_sum_vec10_sink_sel == 75))? _mystream_sum_vec10_sink_wdata : 'hx;
  assign ram_c_10_0_wenable = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                              (_mystream_stream_oready && _mystream_sum_vec10_sink_wenable && (_mystream_sum_vec10_sink_sel == 75))? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_1175;
  assign write_burst_packed_ram_addr_1175 = write_burst_packed_addr_1149 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_1176;
  assign write_burst_packed_ram_wdata_1176 = _myaxi_read_narrow_wdata_1146 >> 352;
  assign ram_c_11_0_wdata = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_wdata_1176 : 
                            (_mystream_stream_oready && _mystream_sum_vec11_sink_wenable && (_mystream_sum_vec11_sink_sel == 76))? _mystream_sum_vec11_sink_wdata : 'hx;
  assign ram_c_11_0_wenable = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                              (_mystream_stream_oready && _mystream_sum_vec11_sink_wenable && (_mystream_sum_vec11_sink_sel == 76))? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_1177;
  assign write_burst_packed_ram_addr_1177 = write_burst_packed_addr_1149 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_1178;
  assign write_burst_packed_ram_wdata_1178 = _myaxi_read_narrow_wdata_1146 >> 384;
  assign ram_c_12_0_wdata = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_wdata_1178 : 
                            (_mystream_stream_oready && _mystream_sum_vec12_sink_wenable && (_mystream_sum_vec12_sink_sel == 77))? _mystream_sum_vec12_sink_wdata : 'hx;
  assign ram_c_12_0_wenable = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                              (_mystream_stream_oready && _mystream_sum_vec12_sink_wenable && (_mystream_sum_vec12_sink_sel == 77))? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_1179;
  assign write_burst_packed_ram_addr_1179 = write_burst_packed_addr_1149 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_1180;
  assign write_burst_packed_ram_wdata_1180 = _myaxi_read_narrow_wdata_1146 >> 416;
  assign ram_c_13_0_wdata = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_wdata_1180 : 
                            (_mystream_stream_oready && _mystream_sum_vec13_sink_wenable && (_mystream_sum_vec13_sink_sel == 78))? _mystream_sum_vec13_sink_wdata : 'hx;
  assign ram_c_13_0_wenable = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                              (_mystream_stream_oready && _mystream_sum_vec13_sink_wenable && (_mystream_sum_vec13_sink_sel == 78))? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_1181;
  assign write_burst_packed_ram_addr_1181 = write_burst_packed_addr_1149 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_1182;
  assign write_burst_packed_ram_wdata_1182 = _myaxi_read_narrow_wdata_1146 >> 448;
  assign ram_c_14_0_wdata = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_wdata_1182 : 
                            (_mystream_stream_oready && _mystream_sum_vec14_sink_wenable && (_mystream_sum_vec14_sink_sel == 79))? _mystream_sum_vec14_sink_wdata : 'hx;
  assign ram_c_14_0_wenable = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                              (_mystream_stream_oready && _mystream_sum_vec14_sink_wenable && (_mystream_sum_vec14_sink_sel == 79))? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_1183;
  assign write_burst_packed_ram_addr_1183 = write_burst_packed_addr_1149 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_1184;
  assign write_burst_packed_ram_wdata_1184 = _myaxi_read_narrow_wdata_1146 >> 480;
  assign ram_c_15_0_wdata = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_wdata_1184 : 
                            (_mystream_stream_oready && _mystream_sum_vec15_sink_wenable && (_mystream_sum_vec15_sink_sel == 80))? _mystream_sum_vec15_sink_wdata : 'hx;
  assign ram_c_15_0_wenable = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                              (_mystream_stream_oready && _mystream_sum_vec15_sink_wenable && (_mystream_sum_vec15_sink_sel == 80))? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_1185;
  assign write_burst_packed_ram_addr_1185 = write_burst_packed_addr_1149 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_1186;
  assign write_burst_packed_ram_wdata_1186 = _myaxi_read_narrow_wdata_1146 >> 512;
  assign ram_c_16_0_wdata = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_wdata_1186 : 
                            (_mystream_stream_oready && _mystream_sum_vec16_sink_wenable && (_mystream_sum_vec16_sink_sel == 81))? _mystream_sum_vec16_sink_wdata : 'hx;
  assign ram_c_16_0_wenable = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                              (_mystream_stream_oready && _mystream_sum_vec16_sink_wenable && (_mystream_sum_vec16_sink_sel == 81))? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_1187;
  assign write_burst_packed_ram_addr_1187 = write_burst_packed_addr_1149 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_1188;
  assign write_burst_packed_ram_wdata_1188 = _myaxi_read_narrow_wdata_1146 >> 544;
  assign ram_c_17_0_wdata = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_wdata_1188 : 
                            (_mystream_stream_oready && _mystream_sum_vec17_sink_wenable && (_mystream_sum_vec17_sink_sel == 82))? _mystream_sum_vec17_sink_wdata : 'hx;
  assign ram_c_17_0_wenable = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                              (_mystream_stream_oready && _mystream_sum_vec17_sink_wenable && (_mystream_sum_vec17_sink_sel == 82))? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_1189;
  assign write_burst_packed_ram_addr_1189 = write_burst_packed_addr_1149 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_1190;
  assign write_burst_packed_ram_wdata_1190 = _myaxi_read_narrow_wdata_1146 >> 576;
  assign ram_c_18_0_wdata = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_wdata_1190 : 
                            (_mystream_stream_oready && _mystream_sum_vec18_sink_wenable && (_mystream_sum_vec18_sink_sel == 83))? _mystream_sum_vec18_sink_wdata : 'hx;
  assign ram_c_18_0_wenable = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                              (_mystream_stream_oready && _mystream_sum_vec18_sink_wenable && (_mystream_sum_vec18_sink_sel == 83))? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_1191;
  assign write_burst_packed_ram_addr_1191 = write_burst_packed_addr_1149 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_1192;
  assign write_burst_packed_ram_wdata_1192 = _myaxi_read_narrow_wdata_1146 >> 608;
  assign ram_c_19_0_wdata = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_wdata_1192 : 
                            (_mystream_stream_oready && _mystream_sum_vec19_sink_wenable && (_mystream_sum_vec19_sink_sel == 84))? _mystream_sum_vec19_sink_wdata : 'hx;
  assign ram_c_19_0_wenable = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                              (_mystream_stream_oready && _mystream_sum_vec19_sink_wenable && (_mystream_sum_vec19_sink_sel == 84))? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_1193;
  assign write_burst_packed_ram_addr_1193 = write_burst_packed_addr_1149 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_1194;
  assign write_burst_packed_ram_wdata_1194 = _myaxi_read_narrow_wdata_1146 >> 640;
  assign ram_c_20_0_wdata = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_wdata_1194 : 
                            (_mystream_stream_oready && _mystream_sum_vec20_sink_wenable && (_mystream_sum_vec20_sink_sel == 85))? _mystream_sum_vec20_sink_wdata : 'hx;
  assign ram_c_20_0_wenable = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                              (_mystream_stream_oready && _mystream_sum_vec20_sink_wenable && (_mystream_sum_vec20_sink_sel == 85))? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_1195;
  assign write_burst_packed_ram_addr_1195 = write_burst_packed_addr_1149 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_1196;
  assign write_burst_packed_ram_wdata_1196 = _myaxi_read_narrow_wdata_1146 >> 672;
  assign ram_c_21_0_wdata = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_wdata_1196 : 
                            (_mystream_stream_oready && _mystream_sum_vec21_sink_wenable && (_mystream_sum_vec21_sink_sel == 86))? _mystream_sum_vec21_sink_wdata : 'hx;
  assign ram_c_21_0_wenable = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                              (_mystream_stream_oready && _mystream_sum_vec21_sink_wenable && (_mystream_sum_vec21_sink_sel == 86))? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_1197;
  assign write_burst_packed_ram_addr_1197 = write_burst_packed_addr_1149 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_1198;
  assign write_burst_packed_ram_wdata_1198 = _myaxi_read_narrow_wdata_1146 >> 704;
  assign ram_c_22_0_wdata = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_wdata_1198 : 
                            (_mystream_stream_oready && _mystream_sum_vec22_sink_wenable && (_mystream_sum_vec22_sink_sel == 87))? _mystream_sum_vec22_sink_wdata : 'hx;
  assign ram_c_22_0_wenable = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                              (_mystream_stream_oready && _mystream_sum_vec22_sink_wenable && (_mystream_sum_vec22_sink_sel == 87))? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_1199;
  assign write_burst_packed_ram_addr_1199 = write_burst_packed_addr_1149 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_1200;
  assign write_burst_packed_ram_wdata_1200 = _myaxi_read_narrow_wdata_1146 >> 736;
  assign ram_c_23_0_wdata = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_wdata_1200 : 
                            (_mystream_stream_oready && _mystream_sum_vec23_sink_wenable && (_mystream_sum_vec23_sink_sel == 88))? _mystream_sum_vec23_sink_wdata : 'hx;
  assign ram_c_23_0_wenable = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                              (_mystream_stream_oready && _mystream_sum_vec23_sink_wenable && (_mystream_sum_vec23_sink_sel == 88))? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_1201;
  assign write_burst_packed_ram_addr_1201 = write_burst_packed_addr_1149 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_1202;
  assign write_burst_packed_ram_wdata_1202 = _myaxi_read_narrow_wdata_1146 >> 768;
  assign ram_c_24_0_wdata = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_wdata_1202 : 
                            (_mystream_stream_oready && _mystream_sum_vec24_sink_wenable && (_mystream_sum_vec24_sink_sel == 89))? _mystream_sum_vec24_sink_wdata : 'hx;
  assign ram_c_24_0_wenable = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                              (_mystream_stream_oready && _mystream_sum_vec24_sink_wenable && (_mystream_sum_vec24_sink_sel == 89))? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_1203;
  assign write_burst_packed_ram_addr_1203 = write_burst_packed_addr_1149 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_1204;
  assign write_burst_packed_ram_wdata_1204 = _myaxi_read_narrow_wdata_1146 >> 800;
  assign ram_c_25_0_wdata = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_wdata_1204 : 
                            (_mystream_stream_oready && _mystream_sum_vec25_sink_wenable && (_mystream_sum_vec25_sink_sel == 90))? _mystream_sum_vec25_sink_wdata : 'hx;
  assign ram_c_25_0_wenable = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                              (_mystream_stream_oready && _mystream_sum_vec25_sink_wenable && (_mystream_sum_vec25_sink_sel == 90))? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_1205;
  assign write_burst_packed_ram_addr_1205 = write_burst_packed_addr_1149 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_1206;
  assign write_burst_packed_ram_wdata_1206 = _myaxi_read_narrow_wdata_1146 >> 832;
  assign ram_c_26_0_wdata = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_wdata_1206 : 
                            (_mystream_stream_oready && _mystream_sum_vec26_sink_wenable && (_mystream_sum_vec26_sink_sel == 91))? _mystream_sum_vec26_sink_wdata : 'hx;
  assign ram_c_26_0_wenable = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                              (_mystream_stream_oready && _mystream_sum_vec26_sink_wenable && (_mystream_sum_vec26_sink_sel == 91))? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_1207;
  assign write_burst_packed_ram_addr_1207 = write_burst_packed_addr_1149 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_1208;
  assign write_burst_packed_ram_wdata_1208 = _myaxi_read_narrow_wdata_1146 >> 864;
  assign ram_c_27_0_wdata = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_wdata_1208 : 
                            (_mystream_stream_oready && _mystream_sum_vec27_sink_wenable && (_mystream_sum_vec27_sink_sel == 92))? _mystream_sum_vec27_sink_wdata : 'hx;
  assign ram_c_27_0_wenable = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                              (_mystream_stream_oready && _mystream_sum_vec27_sink_wenable && (_mystream_sum_vec27_sink_sel == 92))? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_1209;
  assign write_burst_packed_ram_addr_1209 = write_burst_packed_addr_1149 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_1210;
  assign write_burst_packed_ram_wdata_1210 = _myaxi_read_narrow_wdata_1146 >> 896;
  assign ram_c_28_0_wdata = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_wdata_1210 : 
                            (_mystream_stream_oready && _mystream_sum_vec28_sink_wenable && (_mystream_sum_vec28_sink_sel == 93))? _mystream_sum_vec28_sink_wdata : 'hx;
  assign ram_c_28_0_wenable = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                              (_mystream_stream_oready && _mystream_sum_vec28_sink_wenable && (_mystream_sum_vec28_sink_sel == 93))? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_1211;
  assign write_burst_packed_ram_addr_1211 = write_burst_packed_addr_1149 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_1212;
  assign write_burst_packed_ram_wdata_1212 = _myaxi_read_narrow_wdata_1146 >> 928;
  assign ram_c_29_0_wdata = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_wdata_1212 : 
                            (_mystream_stream_oready && _mystream_sum_vec29_sink_wenable && (_mystream_sum_vec29_sink_sel == 94))? _mystream_sum_vec29_sink_wdata : 'hx;
  assign ram_c_29_0_wenable = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                              (_mystream_stream_oready && _mystream_sum_vec29_sink_wenable && (_mystream_sum_vec29_sink_sel == 94))? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_1213;
  assign write_burst_packed_ram_addr_1213 = write_burst_packed_addr_1149 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_1214;
  assign write_burst_packed_ram_wdata_1214 = _myaxi_read_narrow_wdata_1146 >> 960;
  assign ram_c_30_0_wdata = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_wdata_1214 : 
                            (_mystream_stream_oready && _mystream_sum_vec30_sink_wenable && (_mystream_sum_vec30_sink_sel == 95))? _mystream_sum_vec30_sink_wdata : 'hx;
  assign ram_c_30_0_wenable = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                              (_mystream_stream_oready && _mystream_sum_vec30_sink_wenable && (_mystream_sum_vec30_sink_sel == 95))? 1'd1 : 0;
  wire [20-1:0] write_burst_packed_ram_addr_1215;
  assign write_burst_packed_ram_addr_1215 = write_burst_packed_addr_1149 >> 5;
  wire [32-1:0] write_burst_packed_ram_wdata_1216;
  assign write_burst_packed_ram_wdata_1216 = _myaxi_read_narrow_wdata_1146 >> 992;
  assign ram_c_31_0_wdata = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_wdata_1216 : 
                            (_mystream_stream_oready && _mystream_sum_vec31_sink_wenable && (_mystream_sum_vec31_sink_sel == 96))? _mystream_sum_vec31_sink_wdata : 'hx;
  assign ram_c_31_0_wenable = ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                              (_mystream_stream_oready && _mystream_sum_vec31_sink_wenable && (_mystream_sum_vec31_sink_sel == 96))? 1'd1 : 0;
  assign myaxi_rready = (_myaxi_read_data_narrow_fsm == 2) || (_myaxi_read_data_narrow_fsm == 2) || (_myaxi_read_data_fsm == 2) || (_myaxi_read_data_fsm == 2) || (_myaxi_read_data_narrow_fsm == 2);
  reg signed [32-1:0] _th_comp_size_14;
  reg signed [32-1:0] _th_comp_offset_stream_15;
  reg signed [32-1:0] _th_comp_offset_seq_16;
  reg signed [32-1:0] _th_comp_all_ok_17;
  reg signed [32-1:0] _th_comp_i_18;
  wire [5-1:0] read_rtl_bank_1217;
  assign read_rtl_bank_1217 = _th_comp_i_18 + _th_comp_offset_stream_15;
  reg [5-1:0] _tmp_1218;
  localparam _tmp_1219 = 1;
  wire [_tmp_1219-1:0] _tmp_1220;
  assign _tmp_1220 = th_comp == 114;
  reg [_tmp_1219-1:0] __tmp_1220_1;
  localparam _tmp_1221 = 1;
  wire [_tmp_1221-1:0] _tmp_1222;
  assign _tmp_1222 = th_comp == 114;
  reg [_tmp_1221-1:0] __tmp_1222_1;
  localparam _tmp_1223 = 1;
  wire [_tmp_1223-1:0] _tmp_1224;
  assign _tmp_1224 = th_comp == 114;
  reg [_tmp_1223-1:0] __tmp_1224_1;
  localparam _tmp_1225 = 1;
  wire [_tmp_1225-1:0] _tmp_1226;
  assign _tmp_1226 = th_comp == 114;
  reg [_tmp_1225-1:0] __tmp_1226_1;
  localparam _tmp_1227 = 1;
  wire [_tmp_1227-1:0] _tmp_1228;
  assign _tmp_1228 = th_comp == 114;
  reg [_tmp_1227-1:0] __tmp_1228_1;
  localparam _tmp_1229 = 1;
  wire [_tmp_1229-1:0] _tmp_1230;
  assign _tmp_1230 = th_comp == 114;
  reg [_tmp_1229-1:0] __tmp_1230_1;
  localparam _tmp_1231 = 1;
  wire [_tmp_1231-1:0] _tmp_1232;
  assign _tmp_1232 = th_comp == 114;
  reg [_tmp_1231-1:0] __tmp_1232_1;
  localparam _tmp_1233 = 1;
  wire [_tmp_1233-1:0] _tmp_1234;
  assign _tmp_1234 = th_comp == 114;
  reg [_tmp_1233-1:0] __tmp_1234_1;
  localparam _tmp_1235 = 1;
  wire [_tmp_1235-1:0] _tmp_1236;
  assign _tmp_1236 = th_comp == 114;
  reg [_tmp_1235-1:0] __tmp_1236_1;
  localparam _tmp_1237 = 1;
  wire [_tmp_1237-1:0] _tmp_1238;
  assign _tmp_1238 = th_comp == 114;
  reg [_tmp_1237-1:0] __tmp_1238_1;
  localparam _tmp_1239 = 1;
  wire [_tmp_1239-1:0] _tmp_1240;
  assign _tmp_1240 = th_comp == 114;
  reg [_tmp_1239-1:0] __tmp_1240_1;
  localparam _tmp_1241 = 1;
  wire [_tmp_1241-1:0] _tmp_1242;
  assign _tmp_1242 = th_comp == 114;
  reg [_tmp_1241-1:0] __tmp_1242_1;
  localparam _tmp_1243 = 1;
  wire [_tmp_1243-1:0] _tmp_1244;
  assign _tmp_1244 = th_comp == 114;
  reg [_tmp_1243-1:0] __tmp_1244_1;
  localparam _tmp_1245 = 1;
  wire [_tmp_1245-1:0] _tmp_1246;
  assign _tmp_1246 = th_comp == 114;
  reg [_tmp_1245-1:0] __tmp_1246_1;
  localparam _tmp_1247 = 1;
  wire [_tmp_1247-1:0] _tmp_1248;
  assign _tmp_1248 = th_comp == 114;
  reg [_tmp_1247-1:0] __tmp_1248_1;
  localparam _tmp_1249 = 1;
  wire [_tmp_1249-1:0] _tmp_1250;
  assign _tmp_1250 = th_comp == 114;
  reg [_tmp_1249-1:0] __tmp_1250_1;
  localparam _tmp_1251 = 1;
  wire [_tmp_1251-1:0] _tmp_1252;
  assign _tmp_1252 = th_comp == 114;
  reg [_tmp_1251-1:0] __tmp_1252_1;
  localparam _tmp_1253 = 1;
  wire [_tmp_1253-1:0] _tmp_1254;
  assign _tmp_1254 = th_comp == 114;
  reg [_tmp_1253-1:0] __tmp_1254_1;
  localparam _tmp_1255 = 1;
  wire [_tmp_1255-1:0] _tmp_1256;
  assign _tmp_1256 = th_comp == 114;
  reg [_tmp_1255-1:0] __tmp_1256_1;
  localparam _tmp_1257 = 1;
  wire [_tmp_1257-1:0] _tmp_1258;
  assign _tmp_1258 = th_comp == 114;
  reg [_tmp_1257-1:0] __tmp_1258_1;
  localparam _tmp_1259 = 1;
  wire [_tmp_1259-1:0] _tmp_1260;
  assign _tmp_1260 = th_comp == 114;
  reg [_tmp_1259-1:0] __tmp_1260_1;
  localparam _tmp_1261 = 1;
  wire [_tmp_1261-1:0] _tmp_1262;
  assign _tmp_1262 = th_comp == 114;
  reg [_tmp_1261-1:0] __tmp_1262_1;
  localparam _tmp_1263 = 1;
  wire [_tmp_1263-1:0] _tmp_1264;
  assign _tmp_1264 = th_comp == 114;
  reg [_tmp_1263-1:0] __tmp_1264_1;
  localparam _tmp_1265 = 1;
  wire [_tmp_1265-1:0] _tmp_1266;
  assign _tmp_1266 = th_comp == 114;
  reg [_tmp_1265-1:0] __tmp_1266_1;
  localparam _tmp_1267 = 1;
  wire [_tmp_1267-1:0] _tmp_1268;
  assign _tmp_1268 = th_comp == 114;
  reg [_tmp_1267-1:0] __tmp_1268_1;
  localparam _tmp_1269 = 1;
  wire [_tmp_1269-1:0] _tmp_1270;
  assign _tmp_1270 = th_comp == 114;
  reg [_tmp_1269-1:0] __tmp_1270_1;
  localparam _tmp_1271 = 1;
  wire [_tmp_1271-1:0] _tmp_1272;
  assign _tmp_1272 = th_comp == 114;
  reg [_tmp_1271-1:0] __tmp_1272_1;
  localparam _tmp_1273 = 1;
  wire [_tmp_1273-1:0] _tmp_1274;
  assign _tmp_1274 = th_comp == 114;
  reg [_tmp_1273-1:0] __tmp_1274_1;
  localparam _tmp_1275 = 1;
  wire [_tmp_1275-1:0] _tmp_1276;
  assign _tmp_1276 = th_comp == 114;
  reg [_tmp_1275-1:0] __tmp_1276_1;
  localparam _tmp_1277 = 1;
  wire [_tmp_1277-1:0] _tmp_1278;
  assign _tmp_1278 = th_comp == 114;
  reg [_tmp_1277-1:0] __tmp_1278_1;
  localparam _tmp_1279 = 1;
  wire [_tmp_1279-1:0] _tmp_1280;
  assign _tmp_1280 = th_comp == 114;
  reg [_tmp_1279-1:0] __tmp_1280_1;
  localparam _tmp_1281 = 1;
  wire [_tmp_1281-1:0] _tmp_1282;
  assign _tmp_1282 = th_comp == 114;
  reg [_tmp_1281-1:0] __tmp_1282_1;
  wire signed [32-1:0] read_rtl_rdata_1283;
  wire read_rtl_rvalid_1284;
  assign read_rtl_rdata_1283 = (_tmp_1218 == 0)? ram_c_0_0_rdata : 
                               (_tmp_1218 == 1)? ram_c_1_0_rdata : 
                               (_tmp_1218 == 2)? ram_c_2_0_rdata : 
                               (_tmp_1218 == 3)? ram_c_3_0_rdata : 
                               (_tmp_1218 == 4)? ram_c_4_0_rdata : 
                               (_tmp_1218 == 5)? ram_c_5_0_rdata : 
                               (_tmp_1218 == 6)? ram_c_6_0_rdata : 
                               (_tmp_1218 == 7)? ram_c_7_0_rdata : 
                               (_tmp_1218 == 8)? ram_c_8_0_rdata : 
                               (_tmp_1218 == 9)? ram_c_9_0_rdata : 
                               (_tmp_1218 == 10)? ram_c_10_0_rdata : 
                               (_tmp_1218 == 11)? ram_c_11_0_rdata : 
                               (_tmp_1218 == 12)? ram_c_12_0_rdata : 
                               (_tmp_1218 == 13)? ram_c_13_0_rdata : 
                               (_tmp_1218 == 14)? ram_c_14_0_rdata : 
                               (_tmp_1218 == 15)? ram_c_15_0_rdata : 
                               (_tmp_1218 == 16)? ram_c_16_0_rdata : 
                               (_tmp_1218 == 17)? ram_c_17_0_rdata : 
                               (_tmp_1218 == 18)? ram_c_18_0_rdata : 
                               (_tmp_1218 == 19)? ram_c_19_0_rdata : 
                               (_tmp_1218 == 20)? ram_c_20_0_rdata : 
                               (_tmp_1218 == 21)? ram_c_21_0_rdata : 
                               (_tmp_1218 == 22)? ram_c_22_0_rdata : 
                               (_tmp_1218 == 23)? ram_c_23_0_rdata : 
                               (_tmp_1218 == 24)? ram_c_24_0_rdata : 
                               (_tmp_1218 == 25)? ram_c_25_0_rdata : 
                               (_tmp_1218 == 26)? ram_c_26_0_rdata : 
                               (_tmp_1218 == 27)? ram_c_27_0_rdata : 
                               (_tmp_1218 == 28)? ram_c_28_0_rdata : 
                               (_tmp_1218 == 29)? ram_c_29_0_rdata : 
                               (_tmp_1218 == 30)? ram_c_30_0_rdata : 
                               (_tmp_1218 == 31)? ram_c_31_0_rdata : 0;
  assign read_rtl_rvalid_1284 = __tmp_1220_1;
  reg signed [32-1:0] read_rdata_1285;
  reg signed [32-1:0] _th_comp_st_19;
  wire [5-1:0] read_rtl_bank_1286;
  assign read_rtl_bank_1286 = _th_comp_i_18 + _th_comp_offset_seq_16;
  reg [5-1:0] _tmp_1287;
  assign ram_c_0_0_addr = (th_comp == 116)? _th_comp_i_18 + _th_comp_offset_seq_16 >> 5 : 
                          (th_comp == 114)? _th_comp_i_18 + _th_comp_offset_stream_15 >> 5 : 
                          ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_addr_1153 : 
                          (_mystream_stream_oready && _mystream_sum_vec0_sink_wenable && (_mystream_sum_vec0_sink_sel == 65))? _mystream_sum_vec0_sink_waddr : 'hx;
  assign ram_c_0_0_enable = (th_comp == 116)? 1'd1 : 
                            (th_comp == 114)? 1'd1 : 
                            ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                            (_mystream_stream_oready && _mystream_sum_vec0_sink_wenable && (_mystream_sum_vec0_sink_sel == 65))? 1'd1 : 0;
  localparam _tmp_1288 = 1;
  wire [_tmp_1288-1:0] _tmp_1289;
  assign _tmp_1289 = th_comp == 116;
  reg [_tmp_1288-1:0] __tmp_1289_1;
  assign ram_c_1_0_addr = (th_comp == 116)? _th_comp_i_18 + _th_comp_offset_seq_16 >> 5 : 
                          (th_comp == 114)? _th_comp_i_18 + _th_comp_offset_stream_15 >> 5 : 
                          ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_addr_1155 : 
                          (_mystream_stream_oready && _mystream_sum_vec1_sink_wenable && (_mystream_sum_vec1_sink_sel == 66))? _mystream_sum_vec1_sink_waddr : 'hx;
  assign ram_c_1_0_enable = (th_comp == 116)? 1'd1 : 
                            (th_comp == 114)? 1'd1 : 
                            ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                            (_mystream_stream_oready && _mystream_sum_vec1_sink_wenable && (_mystream_sum_vec1_sink_sel == 66))? 1'd1 : 0;
  localparam _tmp_1290 = 1;
  wire [_tmp_1290-1:0] _tmp_1291;
  assign _tmp_1291 = th_comp == 116;
  reg [_tmp_1290-1:0] __tmp_1291_1;
  assign ram_c_2_0_addr = (th_comp == 116)? _th_comp_i_18 + _th_comp_offset_seq_16 >> 5 : 
                          (th_comp == 114)? _th_comp_i_18 + _th_comp_offset_stream_15 >> 5 : 
                          ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_addr_1157 : 
                          (_mystream_stream_oready && _mystream_sum_vec2_sink_wenable && (_mystream_sum_vec2_sink_sel == 67))? _mystream_sum_vec2_sink_waddr : 'hx;
  assign ram_c_2_0_enable = (th_comp == 116)? 1'd1 : 
                            (th_comp == 114)? 1'd1 : 
                            ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                            (_mystream_stream_oready && _mystream_sum_vec2_sink_wenable && (_mystream_sum_vec2_sink_sel == 67))? 1'd1 : 0;
  localparam _tmp_1292 = 1;
  wire [_tmp_1292-1:0] _tmp_1293;
  assign _tmp_1293 = th_comp == 116;
  reg [_tmp_1292-1:0] __tmp_1293_1;
  assign ram_c_3_0_addr = (th_comp == 116)? _th_comp_i_18 + _th_comp_offset_seq_16 >> 5 : 
                          (th_comp == 114)? _th_comp_i_18 + _th_comp_offset_stream_15 >> 5 : 
                          ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_addr_1159 : 
                          (_mystream_stream_oready && _mystream_sum_vec3_sink_wenable && (_mystream_sum_vec3_sink_sel == 68))? _mystream_sum_vec3_sink_waddr : 'hx;
  assign ram_c_3_0_enable = (th_comp == 116)? 1'd1 : 
                            (th_comp == 114)? 1'd1 : 
                            ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                            (_mystream_stream_oready && _mystream_sum_vec3_sink_wenable && (_mystream_sum_vec3_sink_sel == 68))? 1'd1 : 0;
  localparam _tmp_1294 = 1;
  wire [_tmp_1294-1:0] _tmp_1295;
  assign _tmp_1295 = th_comp == 116;
  reg [_tmp_1294-1:0] __tmp_1295_1;
  assign ram_c_4_0_addr = (th_comp == 116)? _th_comp_i_18 + _th_comp_offset_seq_16 >> 5 : 
                          (th_comp == 114)? _th_comp_i_18 + _th_comp_offset_stream_15 >> 5 : 
                          ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_addr_1161 : 
                          (_mystream_stream_oready && _mystream_sum_vec4_sink_wenable && (_mystream_sum_vec4_sink_sel == 69))? _mystream_sum_vec4_sink_waddr : 'hx;
  assign ram_c_4_0_enable = (th_comp == 116)? 1'd1 : 
                            (th_comp == 114)? 1'd1 : 
                            ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                            (_mystream_stream_oready && _mystream_sum_vec4_sink_wenable && (_mystream_sum_vec4_sink_sel == 69))? 1'd1 : 0;
  localparam _tmp_1296 = 1;
  wire [_tmp_1296-1:0] _tmp_1297;
  assign _tmp_1297 = th_comp == 116;
  reg [_tmp_1296-1:0] __tmp_1297_1;
  assign ram_c_5_0_addr = (th_comp == 116)? _th_comp_i_18 + _th_comp_offset_seq_16 >> 5 : 
                          (th_comp == 114)? _th_comp_i_18 + _th_comp_offset_stream_15 >> 5 : 
                          ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_addr_1163 : 
                          (_mystream_stream_oready && _mystream_sum_vec5_sink_wenable && (_mystream_sum_vec5_sink_sel == 70))? _mystream_sum_vec5_sink_waddr : 'hx;
  assign ram_c_5_0_enable = (th_comp == 116)? 1'd1 : 
                            (th_comp == 114)? 1'd1 : 
                            ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                            (_mystream_stream_oready && _mystream_sum_vec5_sink_wenable && (_mystream_sum_vec5_sink_sel == 70))? 1'd1 : 0;
  localparam _tmp_1298 = 1;
  wire [_tmp_1298-1:0] _tmp_1299;
  assign _tmp_1299 = th_comp == 116;
  reg [_tmp_1298-1:0] __tmp_1299_1;
  assign ram_c_6_0_addr = (th_comp == 116)? _th_comp_i_18 + _th_comp_offset_seq_16 >> 5 : 
                          (th_comp == 114)? _th_comp_i_18 + _th_comp_offset_stream_15 >> 5 : 
                          ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_addr_1165 : 
                          (_mystream_stream_oready && _mystream_sum_vec6_sink_wenable && (_mystream_sum_vec6_sink_sel == 71))? _mystream_sum_vec6_sink_waddr : 'hx;
  assign ram_c_6_0_enable = (th_comp == 116)? 1'd1 : 
                            (th_comp == 114)? 1'd1 : 
                            ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                            (_mystream_stream_oready && _mystream_sum_vec6_sink_wenable && (_mystream_sum_vec6_sink_sel == 71))? 1'd1 : 0;
  localparam _tmp_1300 = 1;
  wire [_tmp_1300-1:0] _tmp_1301;
  assign _tmp_1301 = th_comp == 116;
  reg [_tmp_1300-1:0] __tmp_1301_1;
  assign ram_c_7_0_addr = (th_comp == 116)? _th_comp_i_18 + _th_comp_offset_seq_16 >> 5 : 
                          (th_comp == 114)? _th_comp_i_18 + _th_comp_offset_stream_15 >> 5 : 
                          ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_addr_1167 : 
                          (_mystream_stream_oready && _mystream_sum_vec7_sink_wenable && (_mystream_sum_vec7_sink_sel == 72))? _mystream_sum_vec7_sink_waddr : 'hx;
  assign ram_c_7_0_enable = (th_comp == 116)? 1'd1 : 
                            (th_comp == 114)? 1'd1 : 
                            ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                            (_mystream_stream_oready && _mystream_sum_vec7_sink_wenable && (_mystream_sum_vec7_sink_sel == 72))? 1'd1 : 0;
  localparam _tmp_1302 = 1;
  wire [_tmp_1302-1:0] _tmp_1303;
  assign _tmp_1303 = th_comp == 116;
  reg [_tmp_1302-1:0] __tmp_1303_1;
  assign ram_c_8_0_addr = (th_comp == 116)? _th_comp_i_18 + _th_comp_offset_seq_16 >> 5 : 
                          (th_comp == 114)? _th_comp_i_18 + _th_comp_offset_stream_15 >> 5 : 
                          ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_addr_1169 : 
                          (_mystream_stream_oready && _mystream_sum_vec8_sink_wenable && (_mystream_sum_vec8_sink_sel == 73))? _mystream_sum_vec8_sink_waddr : 'hx;
  assign ram_c_8_0_enable = (th_comp == 116)? 1'd1 : 
                            (th_comp == 114)? 1'd1 : 
                            ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                            (_mystream_stream_oready && _mystream_sum_vec8_sink_wenable && (_mystream_sum_vec8_sink_sel == 73))? 1'd1 : 0;
  localparam _tmp_1304 = 1;
  wire [_tmp_1304-1:0] _tmp_1305;
  assign _tmp_1305 = th_comp == 116;
  reg [_tmp_1304-1:0] __tmp_1305_1;
  assign ram_c_9_0_addr = (th_comp == 116)? _th_comp_i_18 + _th_comp_offset_seq_16 >> 5 : 
                          (th_comp == 114)? _th_comp_i_18 + _th_comp_offset_stream_15 >> 5 : 
                          ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_addr_1171 : 
                          (_mystream_stream_oready && _mystream_sum_vec9_sink_wenable && (_mystream_sum_vec9_sink_sel == 74))? _mystream_sum_vec9_sink_waddr : 'hx;
  assign ram_c_9_0_enable = (th_comp == 116)? 1'd1 : 
                            (th_comp == 114)? 1'd1 : 
                            ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                            (_mystream_stream_oready && _mystream_sum_vec9_sink_wenable && (_mystream_sum_vec9_sink_sel == 74))? 1'd1 : 0;
  localparam _tmp_1306 = 1;
  wire [_tmp_1306-1:0] _tmp_1307;
  assign _tmp_1307 = th_comp == 116;
  reg [_tmp_1306-1:0] __tmp_1307_1;
  assign ram_c_10_0_addr = (th_comp == 116)? _th_comp_i_18 + _th_comp_offset_seq_16 >> 5 : 
                           (th_comp == 114)? _th_comp_i_18 + _th_comp_offset_stream_15 >> 5 : 
                           ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_addr_1173 : 
                           (_mystream_stream_oready && _mystream_sum_vec10_sink_wenable && (_mystream_sum_vec10_sink_sel == 75))? _mystream_sum_vec10_sink_waddr : 'hx;
  assign ram_c_10_0_enable = (th_comp == 116)? 1'd1 : 
                             (th_comp == 114)? 1'd1 : 
                             ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                             (_mystream_stream_oready && _mystream_sum_vec10_sink_wenable && (_mystream_sum_vec10_sink_sel == 75))? 1'd1 : 0;
  localparam _tmp_1308 = 1;
  wire [_tmp_1308-1:0] _tmp_1309;
  assign _tmp_1309 = th_comp == 116;
  reg [_tmp_1308-1:0] __tmp_1309_1;
  assign ram_c_11_0_addr = (th_comp == 116)? _th_comp_i_18 + _th_comp_offset_seq_16 >> 5 : 
                           (th_comp == 114)? _th_comp_i_18 + _th_comp_offset_stream_15 >> 5 : 
                           ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_addr_1175 : 
                           (_mystream_stream_oready && _mystream_sum_vec11_sink_wenable && (_mystream_sum_vec11_sink_sel == 76))? _mystream_sum_vec11_sink_waddr : 'hx;
  assign ram_c_11_0_enable = (th_comp == 116)? 1'd1 : 
                             (th_comp == 114)? 1'd1 : 
                             ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                             (_mystream_stream_oready && _mystream_sum_vec11_sink_wenable && (_mystream_sum_vec11_sink_sel == 76))? 1'd1 : 0;
  localparam _tmp_1310 = 1;
  wire [_tmp_1310-1:0] _tmp_1311;
  assign _tmp_1311 = th_comp == 116;
  reg [_tmp_1310-1:0] __tmp_1311_1;
  assign ram_c_12_0_addr = (th_comp == 116)? _th_comp_i_18 + _th_comp_offset_seq_16 >> 5 : 
                           (th_comp == 114)? _th_comp_i_18 + _th_comp_offset_stream_15 >> 5 : 
                           ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_addr_1177 : 
                           (_mystream_stream_oready && _mystream_sum_vec12_sink_wenable && (_mystream_sum_vec12_sink_sel == 77))? _mystream_sum_vec12_sink_waddr : 'hx;
  assign ram_c_12_0_enable = (th_comp == 116)? 1'd1 : 
                             (th_comp == 114)? 1'd1 : 
                             ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                             (_mystream_stream_oready && _mystream_sum_vec12_sink_wenable && (_mystream_sum_vec12_sink_sel == 77))? 1'd1 : 0;
  localparam _tmp_1312 = 1;
  wire [_tmp_1312-1:0] _tmp_1313;
  assign _tmp_1313 = th_comp == 116;
  reg [_tmp_1312-1:0] __tmp_1313_1;
  assign ram_c_13_0_addr = (th_comp == 116)? _th_comp_i_18 + _th_comp_offset_seq_16 >> 5 : 
                           (th_comp == 114)? _th_comp_i_18 + _th_comp_offset_stream_15 >> 5 : 
                           ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_addr_1179 : 
                           (_mystream_stream_oready && _mystream_sum_vec13_sink_wenable && (_mystream_sum_vec13_sink_sel == 78))? _mystream_sum_vec13_sink_waddr : 'hx;
  assign ram_c_13_0_enable = (th_comp == 116)? 1'd1 : 
                             (th_comp == 114)? 1'd1 : 
                             ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                             (_mystream_stream_oready && _mystream_sum_vec13_sink_wenable && (_mystream_sum_vec13_sink_sel == 78))? 1'd1 : 0;
  localparam _tmp_1314 = 1;
  wire [_tmp_1314-1:0] _tmp_1315;
  assign _tmp_1315 = th_comp == 116;
  reg [_tmp_1314-1:0] __tmp_1315_1;
  assign ram_c_14_0_addr = (th_comp == 116)? _th_comp_i_18 + _th_comp_offset_seq_16 >> 5 : 
                           (th_comp == 114)? _th_comp_i_18 + _th_comp_offset_stream_15 >> 5 : 
                           ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_addr_1181 : 
                           (_mystream_stream_oready && _mystream_sum_vec14_sink_wenable && (_mystream_sum_vec14_sink_sel == 79))? _mystream_sum_vec14_sink_waddr : 'hx;
  assign ram_c_14_0_enable = (th_comp == 116)? 1'd1 : 
                             (th_comp == 114)? 1'd1 : 
                             ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                             (_mystream_stream_oready && _mystream_sum_vec14_sink_wenable && (_mystream_sum_vec14_sink_sel == 79))? 1'd1 : 0;
  localparam _tmp_1316 = 1;
  wire [_tmp_1316-1:0] _tmp_1317;
  assign _tmp_1317 = th_comp == 116;
  reg [_tmp_1316-1:0] __tmp_1317_1;
  assign ram_c_15_0_addr = (th_comp == 116)? _th_comp_i_18 + _th_comp_offset_seq_16 >> 5 : 
                           (th_comp == 114)? _th_comp_i_18 + _th_comp_offset_stream_15 >> 5 : 
                           ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_addr_1183 : 
                           (_mystream_stream_oready && _mystream_sum_vec15_sink_wenable && (_mystream_sum_vec15_sink_sel == 80))? _mystream_sum_vec15_sink_waddr : 'hx;
  assign ram_c_15_0_enable = (th_comp == 116)? 1'd1 : 
                             (th_comp == 114)? 1'd1 : 
                             ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                             (_mystream_stream_oready && _mystream_sum_vec15_sink_wenable && (_mystream_sum_vec15_sink_sel == 80))? 1'd1 : 0;
  localparam _tmp_1318 = 1;
  wire [_tmp_1318-1:0] _tmp_1319;
  assign _tmp_1319 = th_comp == 116;
  reg [_tmp_1318-1:0] __tmp_1319_1;
  assign ram_c_16_0_addr = (th_comp == 116)? _th_comp_i_18 + _th_comp_offset_seq_16 >> 5 : 
                           (th_comp == 114)? _th_comp_i_18 + _th_comp_offset_stream_15 >> 5 : 
                           ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_addr_1185 : 
                           (_mystream_stream_oready && _mystream_sum_vec16_sink_wenable && (_mystream_sum_vec16_sink_sel == 81))? _mystream_sum_vec16_sink_waddr : 'hx;
  assign ram_c_16_0_enable = (th_comp == 116)? 1'd1 : 
                             (th_comp == 114)? 1'd1 : 
                             ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                             (_mystream_stream_oready && _mystream_sum_vec16_sink_wenable && (_mystream_sum_vec16_sink_sel == 81))? 1'd1 : 0;
  localparam _tmp_1320 = 1;
  wire [_tmp_1320-1:0] _tmp_1321;
  assign _tmp_1321 = th_comp == 116;
  reg [_tmp_1320-1:0] __tmp_1321_1;
  assign ram_c_17_0_addr = (th_comp == 116)? _th_comp_i_18 + _th_comp_offset_seq_16 >> 5 : 
                           (th_comp == 114)? _th_comp_i_18 + _th_comp_offset_stream_15 >> 5 : 
                           ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_addr_1187 : 
                           (_mystream_stream_oready && _mystream_sum_vec17_sink_wenable && (_mystream_sum_vec17_sink_sel == 82))? _mystream_sum_vec17_sink_waddr : 'hx;
  assign ram_c_17_0_enable = (th_comp == 116)? 1'd1 : 
                             (th_comp == 114)? 1'd1 : 
                             ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                             (_mystream_stream_oready && _mystream_sum_vec17_sink_wenable && (_mystream_sum_vec17_sink_sel == 82))? 1'd1 : 0;
  localparam _tmp_1322 = 1;
  wire [_tmp_1322-1:0] _tmp_1323;
  assign _tmp_1323 = th_comp == 116;
  reg [_tmp_1322-1:0] __tmp_1323_1;
  assign ram_c_18_0_addr = (th_comp == 116)? _th_comp_i_18 + _th_comp_offset_seq_16 >> 5 : 
                           (th_comp == 114)? _th_comp_i_18 + _th_comp_offset_stream_15 >> 5 : 
                           ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_addr_1189 : 
                           (_mystream_stream_oready && _mystream_sum_vec18_sink_wenable && (_mystream_sum_vec18_sink_sel == 83))? _mystream_sum_vec18_sink_waddr : 'hx;
  assign ram_c_18_0_enable = (th_comp == 116)? 1'd1 : 
                             (th_comp == 114)? 1'd1 : 
                             ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                             (_mystream_stream_oready && _mystream_sum_vec18_sink_wenable && (_mystream_sum_vec18_sink_sel == 83))? 1'd1 : 0;
  localparam _tmp_1324 = 1;
  wire [_tmp_1324-1:0] _tmp_1325;
  assign _tmp_1325 = th_comp == 116;
  reg [_tmp_1324-1:0] __tmp_1325_1;
  assign ram_c_19_0_addr = (th_comp == 116)? _th_comp_i_18 + _th_comp_offset_seq_16 >> 5 : 
                           (th_comp == 114)? _th_comp_i_18 + _th_comp_offset_stream_15 >> 5 : 
                           ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_addr_1191 : 
                           (_mystream_stream_oready && _mystream_sum_vec19_sink_wenable && (_mystream_sum_vec19_sink_sel == 84))? _mystream_sum_vec19_sink_waddr : 'hx;
  assign ram_c_19_0_enable = (th_comp == 116)? 1'd1 : 
                             (th_comp == 114)? 1'd1 : 
                             ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                             (_mystream_stream_oready && _mystream_sum_vec19_sink_wenable && (_mystream_sum_vec19_sink_sel == 84))? 1'd1 : 0;
  localparam _tmp_1326 = 1;
  wire [_tmp_1326-1:0] _tmp_1327;
  assign _tmp_1327 = th_comp == 116;
  reg [_tmp_1326-1:0] __tmp_1327_1;
  assign ram_c_20_0_addr = (th_comp == 116)? _th_comp_i_18 + _th_comp_offset_seq_16 >> 5 : 
                           (th_comp == 114)? _th_comp_i_18 + _th_comp_offset_stream_15 >> 5 : 
                           ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_addr_1193 : 
                           (_mystream_stream_oready && _mystream_sum_vec20_sink_wenable && (_mystream_sum_vec20_sink_sel == 85))? _mystream_sum_vec20_sink_waddr : 'hx;
  assign ram_c_20_0_enable = (th_comp == 116)? 1'd1 : 
                             (th_comp == 114)? 1'd1 : 
                             ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                             (_mystream_stream_oready && _mystream_sum_vec20_sink_wenable && (_mystream_sum_vec20_sink_sel == 85))? 1'd1 : 0;
  localparam _tmp_1328 = 1;
  wire [_tmp_1328-1:0] _tmp_1329;
  assign _tmp_1329 = th_comp == 116;
  reg [_tmp_1328-1:0] __tmp_1329_1;
  assign ram_c_21_0_addr = (th_comp == 116)? _th_comp_i_18 + _th_comp_offset_seq_16 >> 5 : 
                           (th_comp == 114)? _th_comp_i_18 + _th_comp_offset_stream_15 >> 5 : 
                           ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_addr_1195 : 
                           (_mystream_stream_oready && _mystream_sum_vec21_sink_wenable && (_mystream_sum_vec21_sink_sel == 86))? _mystream_sum_vec21_sink_waddr : 'hx;
  assign ram_c_21_0_enable = (th_comp == 116)? 1'd1 : 
                             (th_comp == 114)? 1'd1 : 
                             ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                             (_mystream_stream_oready && _mystream_sum_vec21_sink_wenable && (_mystream_sum_vec21_sink_sel == 86))? 1'd1 : 0;
  localparam _tmp_1330 = 1;
  wire [_tmp_1330-1:0] _tmp_1331;
  assign _tmp_1331 = th_comp == 116;
  reg [_tmp_1330-1:0] __tmp_1331_1;
  assign ram_c_22_0_addr = (th_comp == 116)? _th_comp_i_18 + _th_comp_offset_seq_16 >> 5 : 
                           (th_comp == 114)? _th_comp_i_18 + _th_comp_offset_stream_15 >> 5 : 
                           ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_addr_1197 : 
                           (_mystream_stream_oready && _mystream_sum_vec22_sink_wenable && (_mystream_sum_vec22_sink_sel == 87))? _mystream_sum_vec22_sink_waddr : 'hx;
  assign ram_c_22_0_enable = (th_comp == 116)? 1'd1 : 
                             (th_comp == 114)? 1'd1 : 
                             ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                             (_mystream_stream_oready && _mystream_sum_vec22_sink_wenable && (_mystream_sum_vec22_sink_sel == 87))? 1'd1 : 0;
  localparam _tmp_1332 = 1;
  wire [_tmp_1332-1:0] _tmp_1333;
  assign _tmp_1333 = th_comp == 116;
  reg [_tmp_1332-1:0] __tmp_1333_1;
  assign ram_c_23_0_addr = (th_comp == 116)? _th_comp_i_18 + _th_comp_offset_seq_16 >> 5 : 
                           (th_comp == 114)? _th_comp_i_18 + _th_comp_offset_stream_15 >> 5 : 
                           ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_addr_1199 : 
                           (_mystream_stream_oready && _mystream_sum_vec23_sink_wenable && (_mystream_sum_vec23_sink_sel == 88))? _mystream_sum_vec23_sink_waddr : 'hx;
  assign ram_c_23_0_enable = (th_comp == 116)? 1'd1 : 
                             (th_comp == 114)? 1'd1 : 
                             ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                             (_mystream_stream_oready && _mystream_sum_vec23_sink_wenable && (_mystream_sum_vec23_sink_sel == 88))? 1'd1 : 0;
  localparam _tmp_1334 = 1;
  wire [_tmp_1334-1:0] _tmp_1335;
  assign _tmp_1335 = th_comp == 116;
  reg [_tmp_1334-1:0] __tmp_1335_1;
  assign ram_c_24_0_addr = (th_comp == 116)? _th_comp_i_18 + _th_comp_offset_seq_16 >> 5 : 
                           (th_comp == 114)? _th_comp_i_18 + _th_comp_offset_stream_15 >> 5 : 
                           ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_addr_1201 : 
                           (_mystream_stream_oready && _mystream_sum_vec24_sink_wenable && (_mystream_sum_vec24_sink_sel == 89))? _mystream_sum_vec24_sink_waddr : 'hx;
  assign ram_c_24_0_enable = (th_comp == 116)? 1'd1 : 
                             (th_comp == 114)? 1'd1 : 
                             ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                             (_mystream_stream_oready && _mystream_sum_vec24_sink_wenable && (_mystream_sum_vec24_sink_sel == 89))? 1'd1 : 0;
  localparam _tmp_1336 = 1;
  wire [_tmp_1336-1:0] _tmp_1337;
  assign _tmp_1337 = th_comp == 116;
  reg [_tmp_1336-1:0] __tmp_1337_1;
  assign ram_c_25_0_addr = (th_comp == 116)? _th_comp_i_18 + _th_comp_offset_seq_16 >> 5 : 
                           (th_comp == 114)? _th_comp_i_18 + _th_comp_offset_stream_15 >> 5 : 
                           ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_addr_1203 : 
                           (_mystream_stream_oready && _mystream_sum_vec25_sink_wenable && (_mystream_sum_vec25_sink_sel == 90))? _mystream_sum_vec25_sink_waddr : 'hx;
  assign ram_c_25_0_enable = (th_comp == 116)? 1'd1 : 
                             (th_comp == 114)? 1'd1 : 
                             ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                             (_mystream_stream_oready && _mystream_sum_vec25_sink_wenable && (_mystream_sum_vec25_sink_sel == 90))? 1'd1 : 0;
  localparam _tmp_1338 = 1;
  wire [_tmp_1338-1:0] _tmp_1339;
  assign _tmp_1339 = th_comp == 116;
  reg [_tmp_1338-1:0] __tmp_1339_1;
  assign ram_c_26_0_addr = (th_comp == 116)? _th_comp_i_18 + _th_comp_offset_seq_16 >> 5 : 
                           (th_comp == 114)? _th_comp_i_18 + _th_comp_offset_stream_15 >> 5 : 
                           ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_addr_1205 : 
                           (_mystream_stream_oready && _mystream_sum_vec26_sink_wenable && (_mystream_sum_vec26_sink_sel == 91))? _mystream_sum_vec26_sink_waddr : 'hx;
  assign ram_c_26_0_enable = (th_comp == 116)? 1'd1 : 
                             (th_comp == 114)? 1'd1 : 
                             ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                             (_mystream_stream_oready && _mystream_sum_vec26_sink_wenable && (_mystream_sum_vec26_sink_sel == 91))? 1'd1 : 0;
  localparam _tmp_1340 = 1;
  wire [_tmp_1340-1:0] _tmp_1341;
  assign _tmp_1341 = th_comp == 116;
  reg [_tmp_1340-1:0] __tmp_1341_1;
  assign ram_c_27_0_addr = (th_comp == 116)? _th_comp_i_18 + _th_comp_offset_seq_16 >> 5 : 
                           (th_comp == 114)? _th_comp_i_18 + _th_comp_offset_stream_15 >> 5 : 
                           ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_addr_1207 : 
                           (_mystream_stream_oready && _mystream_sum_vec27_sink_wenable && (_mystream_sum_vec27_sink_sel == 92))? _mystream_sum_vec27_sink_waddr : 'hx;
  assign ram_c_27_0_enable = (th_comp == 116)? 1'd1 : 
                             (th_comp == 114)? 1'd1 : 
                             ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                             (_mystream_stream_oready && _mystream_sum_vec27_sink_wenable && (_mystream_sum_vec27_sink_sel == 92))? 1'd1 : 0;
  localparam _tmp_1342 = 1;
  wire [_tmp_1342-1:0] _tmp_1343;
  assign _tmp_1343 = th_comp == 116;
  reg [_tmp_1342-1:0] __tmp_1343_1;
  assign ram_c_28_0_addr = (th_comp == 116)? _th_comp_i_18 + _th_comp_offset_seq_16 >> 5 : 
                           (th_comp == 114)? _th_comp_i_18 + _th_comp_offset_stream_15 >> 5 : 
                           ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_addr_1209 : 
                           (_mystream_stream_oready && _mystream_sum_vec28_sink_wenable && (_mystream_sum_vec28_sink_sel == 93))? _mystream_sum_vec28_sink_waddr : 'hx;
  assign ram_c_28_0_enable = (th_comp == 116)? 1'd1 : 
                             (th_comp == 114)? 1'd1 : 
                             ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                             (_mystream_stream_oready && _mystream_sum_vec28_sink_wenable && (_mystream_sum_vec28_sink_sel == 93))? 1'd1 : 0;
  localparam _tmp_1344 = 1;
  wire [_tmp_1344-1:0] _tmp_1345;
  assign _tmp_1345 = th_comp == 116;
  reg [_tmp_1344-1:0] __tmp_1345_1;
  assign ram_c_29_0_addr = (th_comp == 116)? _th_comp_i_18 + _th_comp_offset_seq_16 >> 5 : 
                           (th_comp == 114)? _th_comp_i_18 + _th_comp_offset_stream_15 >> 5 : 
                           ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_addr_1211 : 
                           (_mystream_stream_oready && _mystream_sum_vec29_sink_wenable && (_mystream_sum_vec29_sink_sel == 94))? _mystream_sum_vec29_sink_waddr : 'hx;
  assign ram_c_29_0_enable = (th_comp == 116)? 1'd1 : 
                             (th_comp == 114)? 1'd1 : 
                             ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                             (_mystream_stream_oready && _mystream_sum_vec29_sink_wenable && (_mystream_sum_vec29_sink_sel == 94))? 1'd1 : 0;
  localparam _tmp_1346 = 1;
  wire [_tmp_1346-1:0] _tmp_1347;
  assign _tmp_1347 = th_comp == 116;
  reg [_tmp_1346-1:0] __tmp_1347_1;
  assign ram_c_30_0_addr = (th_comp == 116)? _th_comp_i_18 + _th_comp_offset_seq_16 >> 5 : 
                           (th_comp == 114)? _th_comp_i_18 + _th_comp_offset_stream_15 >> 5 : 
                           ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_addr_1213 : 
                           (_mystream_stream_oready && _mystream_sum_vec30_sink_wenable && (_mystream_sum_vec30_sink_sel == 95))? _mystream_sum_vec30_sink_waddr : 'hx;
  assign ram_c_30_0_enable = (th_comp == 116)? 1'd1 : 
                             (th_comp == 114)? 1'd1 : 
                             ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                             (_mystream_stream_oready && _mystream_sum_vec30_sink_wenable && (_mystream_sum_vec30_sink_sel == 95))? 1'd1 : 0;
  localparam _tmp_1348 = 1;
  wire [_tmp_1348-1:0] _tmp_1349;
  assign _tmp_1349 = th_comp == 116;
  reg [_tmp_1348-1:0] __tmp_1349_1;
  assign ram_c_31_0_addr = (th_comp == 116)? _th_comp_i_18 + _th_comp_offset_seq_16 >> 5 : 
                           (th_comp == 114)? _th_comp_i_18 + _th_comp_offset_stream_15 >> 5 : 
                           ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? write_burst_packed_ram_addr_1215 : 
                           (_mystream_stream_oready && _mystream_sum_vec31_sink_wenable && (_mystream_sum_vec31_sink_sel == 96))? _mystream_sum_vec31_sink_waddr : 'hx;
  assign ram_c_31_0_enable = (th_comp == 116)? 1'd1 : 
                             (th_comp == 114)? 1'd1 : 
                             ((write_burst_packed_fsm_5 == 1) && _myaxi_read_narrow_wvalid_1147)? 1'd1 : 
                             (_mystream_stream_oready && _mystream_sum_vec31_sink_wenable && (_mystream_sum_vec31_sink_sel == 96))? 1'd1 : 0;
  localparam _tmp_1350 = 1;
  wire [_tmp_1350-1:0] _tmp_1351;
  assign _tmp_1351 = th_comp == 116;
  reg [_tmp_1350-1:0] __tmp_1351_1;
  wire signed [32-1:0] read_rtl_rdata_1352;
  wire read_rtl_rvalid_1353;
  assign read_rtl_rdata_1352 = (_tmp_1287 == 0)? ram_c_0_0_rdata : 
                               (_tmp_1287 == 1)? ram_c_1_0_rdata : 
                               (_tmp_1287 == 2)? ram_c_2_0_rdata : 
                               (_tmp_1287 == 3)? ram_c_3_0_rdata : 
                               (_tmp_1287 == 4)? ram_c_4_0_rdata : 
                               (_tmp_1287 == 5)? ram_c_5_0_rdata : 
                               (_tmp_1287 == 6)? ram_c_6_0_rdata : 
                               (_tmp_1287 == 7)? ram_c_7_0_rdata : 
                               (_tmp_1287 == 8)? ram_c_8_0_rdata : 
                               (_tmp_1287 == 9)? ram_c_9_0_rdata : 
                               (_tmp_1287 == 10)? ram_c_10_0_rdata : 
                               (_tmp_1287 == 11)? ram_c_11_0_rdata : 
                               (_tmp_1287 == 12)? ram_c_12_0_rdata : 
                               (_tmp_1287 == 13)? ram_c_13_0_rdata : 
                               (_tmp_1287 == 14)? ram_c_14_0_rdata : 
                               (_tmp_1287 == 15)? ram_c_15_0_rdata : 
                               (_tmp_1287 == 16)? ram_c_16_0_rdata : 
                               (_tmp_1287 == 17)? ram_c_17_0_rdata : 
                               (_tmp_1287 == 18)? ram_c_18_0_rdata : 
                               (_tmp_1287 == 19)? ram_c_19_0_rdata : 
                               (_tmp_1287 == 20)? ram_c_20_0_rdata : 
                               (_tmp_1287 == 21)? ram_c_21_0_rdata : 
                               (_tmp_1287 == 22)? ram_c_22_0_rdata : 
                               (_tmp_1287 == 23)? ram_c_23_0_rdata : 
                               (_tmp_1287 == 24)? ram_c_24_0_rdata : 
                               (_tmp_1287 == 25)? ram_c_25_0_rdata : 
                               (_tmp_1287 == 26)? ram_c_26_0_rdata : 
                               (_tmp_1287 == 27)? ram_c_27_0_rdata : 
                               (_tmp_1287 == 28)? ram_c_28_0_rdata : 
                               (_tmp_1287 == 29)? ram_c_29_0_rdata : 
                               (_tmp_1287 == 30)? ram_c_30_0_rdata : 
                               (_tmp_1287 == 31)? ram_c_31_0_rdata : 0;
  assign read_rtl_rvalid_1353 = __tmp_1289_1;
  reg signed [32-1:0] read_rdata_1354;
  reg signed [32-1:0] _th_comp_sq_20;

  always @(posedge CLK) begin
    if(RST) begin
      outstanding_wcount_0 <= 0;
      _myaxi_read_start <= 0;
      _myaxi_write_start <= 0;
      _myaxi_read_op_sel <= 0;
      _myaxi_read_global_addr <= 0;
      _myaxi_read_global_size <= 0;
      _myaxi_read_local_addr <= 0;
      _myaxi_read_local_stride <= 0;
      _myaxi_read_local_size <= 0;
      _myaxi_read_local_blocksize <= 0;
      _myaxi_read_req_idle <= 1;
      _myaxi_read_cur_global_size <= 0;
      myaxi_araddr <= 0;
      myaxi_arlen <= 0;
      myaxi_arvalid <= 0;
      _myaxi_cond_0_1 <= 0;
      _myaxi_read_data_idle <= 1;
      _myaxi_read_op_sel_buf <= 0;
      _myaxi_read_local_addr_buf <= 0;
      _myaxi_read_local_stride_buf <= 0;
      _myaxi_read_local_size_buf <= 0;
      _myaxi_read_local_blocksize_buf <= 0;
      _myaxi_write_op_sel <= 0;
      _myaxi_write_global_addr <= 0;
      _myaxi_write_global_size <= 0;
      _myaxi_write_local_addr <= 0;
      _myaxi_write_local_stride <= 0;
      _myaxi_write_local_size <= 0;
      _myaxi_write_local_blocksize <= 0;
      _myaxi_write_req_idle <= 1;
      _myaxi_write_cur_global_size <= 0;
      myaxi_awaddr <= 0;
      myaxi_awlen <= 0;
      myaxi_awvalid <= 0;
      _myaxi_cond_1_1 <= 0;
      _myaxi_write_data_idle <= 1;
      _myaxi_write_op_sel_buf <= 0;
      _myaxi_write_local_addr_buf <= 0;
      _myaxi_write_local_stride_buf <= 0;
      _myaxi_write_size_buf <= 0;
      _myaxi_write_local_blocksize_buf <= 0;
      myaxi_wdata <= 0;
      myaxi_wvalid <= 0;
      myaxi_wlast <= 0;
      myaxi_wstrb <= 0;
      _myaxi_cond_2_1 <= 0;
    end else begin
      if(_myaxi_cond_0_1) begin
        myaxi_arvalid <= 0;
      end 
      if(_myaxi_cond_1_1) begin
        myaxi_awvalid <= 0;
      end 
      if(_myaxi_cond_2_1) begin
        myaxi_wvalid <= 0;
        myaxi_wlast <= 0;
      end 
      if(myaxi_awvalid && myaxi_awready && !(myaxi_bvalid && myaxi_bready) && (outstanding_wcount_0 < 7)) begin
        outstanding_wcount_0 <= outstanding_wcount_0 + 1;
      end 
      if(!(myaxi_awvalid && myaxi_awready) && (myaxi_bvalid && myaxi_bready) && (outstanding_wcount_0 > 0)) begin
        outstanding_wcount_0 <= outstanding_wcount_0 - 1;
      end 
      _myaxi_read_start <= 0;
      _myaxi_write_start <= 0;
      if((th_comp == 4) && _myaxi_read_req_idle) begin
        _myaxi_read_start <= 1;
        _myaxi_read_op_sel <= 1;
        _myaxi_read_global_addr <= mask_addr_masked_15;
        _myaxi_read_global_size <= _dma_read_packed_local_packed_size_13 << 5;
        _myaxi_read_local_addr <= _th_comp_offset_2;
        _myaxi_read_local_stride <= 32;
        _myaxi_read_local_size <= _dma_read_packed_local_packed_size_13;
        _myaxi_read_local_blocksize <= 1;
      end 
      if((_myaxi_read_req_fsm == 0) && _myaxi_read_start) begin
        _myaxi_read_req_idle <= 0;
      end 
      if(_myaxi_read_start && _myaxi_read_req_fifo_almost_full) begin
        _myaxi_read_start <= 1;
      end 
      if((_myaxi_read_req_fsm == 0) && (_myaxi_read_start || _myaxi_read_cont) && !_myaxi_read_req_fifo_almost_full && (_myaxi_read_global_size <= 256) && ((mask_addr_masked_25 & 4095) + (_myaxi_read_global_size << 2) >= 4096)) begin
        _myaxi_read_cur_global_size <= 4096 - (mask_addr_masked_27 & 4095) >> 2;
        _myaxi_read_global_size <= _myaxi_read_global_size - (4096 - (mask_addr_masked_29 & 4095) >> 2);
      end else if((_myaxi_read_req_fsm == 0) && (_myaxi_read_start || _myaxi_read_cont) && !_myaxi_read_req_fifo_almost_full && (_myaxi_read_global_size <= 256)) begin
        _myaxi_read_cur_global_size <= _myaxi_read_global_size;
        _myaxi_read_global_size <= 0;
      end else if((_myaxi_read_req_fsm == 0) && (_myaxi_read_start || _myaxi_read_cont) && !_myaxi_read_req_fifo_almost_full && ((mask_addr_masked_31 & 4095) + 1024 >= 4096)) begin
        _myaxi_read_cur_global_size <= 4096 - (mask_addr_masked_33 & 4095) >> 2;
        _myaxi_read_global_size <= _myaxi_read_global_size - (4096 - (mask_addr_masked_35 & 4095) >> 2);
      end else if((_myaxi_read_req_fsm == 0) && (_myaxi_read_start || _myaxi_read_cont) && !_myaxi_read_req_fifo_almost_full) begin
        _myaxi_read_cur_global_size <= 256;
        _myaxi_read_global_size <= _myaxi_read_global_size - 256;
      end 
      if((_myaxi_read_req_fsm == 1) && (myaxi_arready || !myaxi_arvalid)) begin
        myaxi_araddr <= _myaxi_read_global_addr;
        myaxi_arlen <= _myaxi_read_cur_global_size - 1;
        myaxi_arvalid <= 1;
      end 
      _myaxi_cond_0_1 <= 1;
      if(myaxi_arvalid && !myaxi_arready) begin
        myaxi_arvalid <= myaxi_arvalid;
      end 
      if((_myaxi_read_req_fsm == 1) && (myaxi_arready || !myaxi_arvalid)) begin
        _myaxi_read_global_addr <= _myaxi_read_global_addr + (_myaxi_read_cur_global_size << 2);
      end 
      if((_myaxi_read_req_fsm == 1) && (myaxi_arready || !myaxi_arvalid) && (_myaxi_read_global_size == 0)) begin
        _myaxi_read_req_idle <= 1;
      end 
      if((_myaxi_read_data_narrow_fsm == 0) && (_myaxi_read_data_idle && !_myaxi_read_req_fifo_empty && (_myaxi_read_op_sel_fifo == 1))) begin
        _myaxi_read_data_idle <= 0;
        _myaxi_read_op_sel_buf <= _myaxi_read_op_sel_fifo;
        _myaxi_read_local_addr_buf <= _myaxi_read_local_addr_fifo;
        _myaxi_read_local_stride_buf <= _myaxi_read_local_stride_fifo;
        _myaxi_read_local_size_buf <= _myaxi_read_local_size_fifo;
        _myaxi_read_local_blocksize_buf <= _myaxi_read_local_blocksize_fifo;
      end 
      if((_myaxi_read_data_narrow_fsm == 2) && (_myaxi_read_op_sel_buf == 1) && myaxi_rvalid && (_myaxi_read_narrow_count_38 == 31)) begin
        _myaxi_read_local_size_buf <= _myaxi_read_local_size_buf - 1;
      end 
      if((_myaxi_read_data_narrow_fsm == 2) && (_myaxi_read_op_sel_buf == 1) && myaxi_rvalid && (_myaxi_read_local_size_buf <= 1) && (_myaxi_read_narrow_count_38 == 31)) begin
        _myaxi_read_data_idle <= 1;
      end 
      if((th_comp == 6) && _myaxi_read_req_idle) begin
        _myaxi_read_start <= 1;
        _myaxi_read_op_sel <= 2;
        _myaxi_read_global_addr <= mask_addr_masked_111;
        _myaxi_read_global_size <= _dma_read_packed_local_packed_size_109 << 5;
        _myaxi_read_local_addr <= _th_comp_offset_2;
        _myaxi_read_local_stride <= 32;
        _myaxi_read_local_size <= _dma_read_packed_local_packed_size_109;
        _myaxi_read_local_blocksize <= 1;
      end 
      if((_myaxi_read_data_narrow_fsm == 0) && (_myaxi_read_data_idle && !_myaxi_read_req_fifo_empty && (_myaxi_read_op_sel_fifo == 2))) begin
        _myaxi_read_data_idle <= 0;
        _myaxi_read_op_sel_buf <= _myaxi_read_op_sel_fifo;
        _myaxi_read_local_addr_buf <= _myaxi_read_local_addr_fifo;
        _myaxi_read_local_stride_buf <= _myaxi_read_local_stride_fifo;
        _myaxi_read_local_size_buf <= _myaxi_read_local_size_fifo;
        _myaxi_read_local_blocksize_buf <= _myaxi_read_local_blocksize_fifo;
      end 
      if((_myaxi_read_data_narrow_fsm == 2) && (_myaxi_read_op_sel_buf == 2) && myaxi_rvalid && (_myaxi_read_narrow_count_114 == 31)) begin
        _myaxi_read_local_size_buf <= _myaxi_read_local_size_buf - 1;
      end 
      if((_myaxi_read_data_narrow_fsm == 2) && (_myaxi_read_op_sel_buf == 2) && myaxi_rvalid && (_myaxi_read_local_size_buf <= 1) && (_myaxi_read_narrow_count_114 == 31)) begin
        _myaxi_read_data_idle <= 1;
      end 
      if((th_comp == 91) && _myaxi_read_req_idle) begin
        _myaxi_read_start <= 1;
        _myaxi_read_op_sel <= 3;
        _myaxi_read_global_addr <= mask_addr_masked_1086;
        _myaxi_read_global_size <= _th_comp_size_0;
        _myaxi_read_local_addr <= _th_comp_offset_2;
        _myaxi_read_local_stride <= 1;
        _myaxi_read_local_size <= _th_comp_size_0;
        _myaxi_read_local_blocksize <= 1;
      end 
      if((_myaxi_read_data_fsm == 0) && (_myaxi_read_data_idle && !_myaxi_read_req_fifo_empty && (_myaxi_read_op_sel_fifo == 3))) begin
        _myaxi_read_data_idle <= 0;
        _myaxi_read_op_sel_buf <= _myaxi_read_op_sel_fifo;
        _myaxi_read_local_addr_buf <= _myaxi_read_local_addr_fifo;
        _myaxi_read_local_stride_buf <= _myaxi_read_local_stride_fifo;
        _myaxi_read_local_size_buf <= _myaxi_read_local_size_fifo;
        _myaxi_read_local_blocksize_buf <= _myaxi_read_local_blocksize_fifo;
      end 
      if((_myaxi_read_data_fsm == 2) && myaxi_rvalid) begin
        _myaxi_read_local_size_buf <= _myaxi_read_local_size_buf - 1;
      end 
      if((_myaxi_read_data_fsm == 2) && myaxi_rvalid && (_myaxi_read_local_size_buf <= 1)) begin
        _myaxi_read_data_idle <= 1;
      end 
      if((th_comp == 93) && _myaxi_read_req_idle) begin
        _myaxi_read_start <= 1;
        _myaxi_read_op_sel <= 4;
        _myaxi_read_global_addr <= mask_addr_masked_1092;
        _myaxi_read_global_size <= _th_comp_size_0;
        _myaxi_read_local_addr <= _th_comp_offset_2;
        _myaxi_read_local_stride <= 1;
        _myaxi_read_local_size <= _th_comp_size_0;
        _myaxi_read_local_blocksize <= 1;
      end 
      if((_myaxi_read_data_fsm == 0) && (_myaxi_read_data_idle && !_myaxi_read_req_fifo_empty && (_myaxi_read_op_sel_fifo == 4))) begin
        _myaxi_read_data_idle <= 0;
        _myaxi_read_op_sel_buf <= _myaxi_read_op_sel_fifo;
        _myaxi_read_local_addr_buf <= _myaxi_read_local_addr_fifo;
        _myaxi_read_local_stride_buf <= _myaxi_read_local_stride_fifo;
        _myaxi_read_local_size_buf <= _myaxi_read_local_size_fifo;
        _myaxi_read_local_blocksize_buf <= _myaxi_read_local_blocksize_fifo;
      end 
      if((_myaxi_read_data_fsm == 2) && myaxi_rvalid) begin
        _myaxi_read_local_size_buf <= _myaxi_read_local_size_buf - 1;
      end 
      if((_myaxi_read_data_fsm == 2) && myaxi_rvalid && (_myaxi_read_local_size_buf <= 1)) begin
        _myaxi_read_data_idle <= 1;
      end 
      if((th_comp == 106) && _myaxi_write_req_idle) begin
        _myaxi_write_start <= 1;
        _myaxi_write_op_sel <= 1;
        _myaxi_write_global_addr <= mask_addr_masked_1104;
        _myaxi_write_global_size <= _th_comp_size_0;
        _myaxi_write_local_addr <= _th_comp_offset_2;
        _myaxi_write_local_stride <= 1;
        _myaxi_write_local_size <= _th_comp_size_0;
        _myaxi_write_local_blocksize <= 1;
      end 
      if((_myaxi_write_req_fsm == 0) && _myaxi_write_start) begin
        _myaxi_write_req_idle <= 0;
      end 
      if(_myaxi_write_start && _myaxi_write_req_fifo_almost_full) begin
        _myaxi_write_start <= 1;
      end 
      if((_myaxi_write_req_fsm == 0) && (_myaxi_write_start || _myaxi_write_cont) && !_myaxi_write_req_fifo_almost_full && (_myaxi_write_global_size <= 256) && ((mask_addr_masked_1114 & 4095) + (_myaxi_write_global_size << 2) >= 4096)) begin
        _myaxi_write_cur_global_size <= 4096 - (mask_addr_masked_1116 & 4095) >> 2;
        _myaxi_write_global_size <= _myaxi_write_global_size - (4096 - (mask_addr_masked_1118 & 4095) >> 2);
      end else if((_myaxi_write_req_fsm == 0) && (_myaxi_write_start || _myaxi_write_cont) && !_myaxi_write_req_fifo_almost_full && (_myaxi_write_global_size <= 256)) begin
        _myaxi_write_cur_global_size <= _myaxi_write_global_size;
        _myaxi_write_global_size <= 0;
      end else if((_myaxi_write_req_fsm == 0) && (_myaxi_write_start || _myaxi_write_cont) && !_myaxi_write_req_fifo_almost_full && ((mask_addr_masked_1120 & 4095) + 1024 >= 4096)) begin
        _myaxi_write_cur_global_size <= 4096 - (mask_addr_masked_1122 & 4095) >> 2;
        _myaxi_write_global_size <= _myaxi_write_global_size - (4096 - (mask_addr_masked_1124 & 4095) >> 2);
      end else if((_myaxi_write_req_fsm == 0) && (_myaxi_write_start || _myaxi_write_cont) && !_myaxi_write_req_fifo_almost_full) begin
        _myaxi_write_cur_global_size <= 256;
        _myaxi_write_global_size <= _myaxi_write_global_size - 256;
      end 
      if((_myaxi_write_req_fsm == 1) && !_myaxi_write_req_fifo_almost_full && (outstanding_wcount_0 < 6) && ((outstanding_wcount_0 < 6) && (myaxi_awready || !myaxi_awvalid))) begin
        myaxi_awaddr <= _myaxi_write_global_addr;
        myaxi_awlen <= _myaxi_write_cur_global_size - 1;
        myaxi_awvalid <= 1;
      end 
      if((_myaxi_write_req_fsm == 1) && !_myaxi_write_req_fifo_almost_full && (outstanding_wcount_0 < 6) && ((outstanding_wcount_0 < 6) && (myaxi_awready || !myaxi_awvalid)) && (_myaxi_write_cur_global_size == 0)) begin
        myaxi_awvalid <= 0;
      end 
      _myaxi_cond_1_1 <= 1;
      if(myaxi_awvalid && !myaxi_awready) begin
        myaxi_awvalid <= myaxi_awvalid;
      end 
      if((_myaxi_write_req_fsm == 1) && ((_myaxi_write_req_fsm == 1) && !_myaxi_write_req_fifo_almost_full && (myaxi_awready || !myaxi_awvalid) && (outstanding_wcount_0 < 6))) begin
        _myaxi_write_global_addr <= _myaxi_write_global_addr + (_myaxi_write_cur_global_size << 2);
      end 
      if((_myaxi_write_req_fsm == 1) && ((_myaxi_write_req_fsm == 1) && !_myaxi_write_req_fifo_almost_full && (myaxi_awready || !myaxi_awvalid) && (outstanding_wcount_0 < 6)) && (_myaxi_write_global_size == 0)) begin
        _myaxi_write_req_idle <= 1;
      end 
      if((_myaxi_write_data_fsm == 0) && (_myaxi_write_data_idle && !_myaxi_write_req_fifo_empty && (_myaxi_write_op_sel_fifo == 1))) begin
        _myaxi_write_data_idle <= 0;
        _myaxi_write_op_sel_buf <= _myaxi_write_op_sel_fifo;
        _myaxi_write_local_addr_buf <= _myaxi_write_local_addr_fifo;
        _myaxi_write_local_stride_buf <= _myaxi_write_local_stride_fifo;
        _myaxi_write_size_buf <= _myaxi_write_size_fifo;
        _myaxi_write_local_blocksize_buf <= _myaxi_write_local_blocksize_fifo;
      end 
      if(_myaxi_write_data_fsm == 1) begin
        _myaxi_write_size_buf <= 0;
      end 
      if((_myaxi_write_data_fsm == 2) && (!_myaxi_write_req_fifo_empty && (_myaxi_write_size_buf == 0))) begin
        _myaxi_write_size_buf <= _myaxi_write_size_fifo;
      end 
      if((_myaxi_write_op_sel_buf == 1) && read_burst_rvalid_1136 && ((myaxi_wready || !myaxi_wvalid) && (_myaxi_write_size_buf > 0)) && (myaxi_wready || !myaxi_wvalid)) begin
        myaxi_wdata <= read_burst_rdata_1140;
        myaxi_wvalid <= 1;
        myaxi_wlast <= read_burst_rlast_1137 || (_myaxi_write_size_buf == 1);
        myaxi_wstrb <= { 4{ 1'd1 } };
      end 
      _myaxi_cond_2_1 <= 1;
      if(myaxi_wvalid && !myaxi_wready) begin
        myaxi_wvalid <= myaxi_wvalid;
        myaxi_wlast <= myaxi_wlast;
      end 
      if((_myaxi_write_data_fsm == 2) && read_burst_rvalid_1136 && ((myaxi_wready || !myaxi_wvalid) && (_myaxi_write_size_buf > 0))) begin
        _myaxi_write_size_buf <= _myaxi_write_size_buf - 1;
      end 
      if((_myaxi_write_data_fsm == 2) && ((_myaxi_write_op_sel_buf == 1) && read_burst_rvalid_1136 && ((myaxi_wready || !myaxi_wvalid) && (_myaxi_write_size_buf > 0))) && read_burst_rlast_1137) begin
        _myaxi_write_data_idle <= 1;
      end 
      if((th_comp == 108) && _myaxi_read_req_idle) begin
        _myaxi_read_start <= 1;
        _myaxi_read_op_sel <= 5;
        _myaxi_read_global_addr <= mask_addr_masked_1145;
        _myaxi_read_global_size <= _dma_read_packed_local_packed_size_1143 << 5;
        _myaxi_read_local_addr <= _th_comp_offset_2;
        _myaxi_read_local_stride <= 32;
        _myaxi_read_local_size <= _dma_read_packed_local_packed_size_1143;
        _myaxi_read_local_blocksize <= 1;
      end 
      if((_myaxi_read_data_narrow_fsm == 0) && (_myaxi_read_data_idle && !_myaxi_read_req_fifo_empty && (_myaxi_read_op_sel_fifo == 5))) begin
        _myaxi_read_data_idle <= 0;
        _myaxi_read_op_sel_buf <= _myaxi_read_op_sel_fifo;
        _myaxi_read_local_addr_buf <= _myaxi_read_local_addr_fifo;
        _myaxi_read_local_stride_buf <= _myaxi_read_local_stride_fifo;
        _myaxi_read_local_size_buf <= _myaxi_read_local_size_fifo;
        _myaxi_read_local_blocksize_buf <= _myaxi_read_local_blocksize_fifo;
      end 
      if((_myaxi_read_data_narrow_fsm == 2) && (_myaxi_read_op_sel_buf == 5) && myaxi_rvalid && (_myaxi_read_narrow_count_1148 == 31)) begin
        _myaxi_read_local_size_buf <= _myaxi_read_local_size_buf - 1;
      end 
      if((_myaxi_read_data_narrow_fsm == 2) && (_myaxi_read_op_sel_buf == 5) && myaxi_rvalid && (_myaxi_read_local_size_buf <= 1) && (_myaxi_read_narrow_count_1148 == 31)) begin
        _myaxi_read_data_idle <= 1;
      end 
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      count__myaxi_read_req_fifo <= 0;
      __tmp_23_1 <= 0;
    end else begin
      if(_myaxi_read_req_fifo_enq && !_myaxi_read_req_fifo_full && (_myaxi_read_req_fifo_deq && !_myaxi_read_req_fifo_empty)) begin
        count__myaxi_read_req_fifo <= count__myaxi_read_req_fifo;
      end else if(_myaxi_read_req_fifo_enq && !_myaxi_read_req_fifo_full) begin
        count__myaxi_read_req_fifo <= count__myaxi_read_req_fifo + 1;
      end else if(_myaxi_read_req_fifo_deq && !_myaxi_read_req_fifo_empty) begin
        count__myaxi_read_req_fifo <= count__myaxi_read_req_fifo - 1;
      end 
      __tmp_23_1 <= _tmp_23;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      count__myaxi_write_req_fifo <= 0;
      __tmp_1112_1 <= 0;
      __tmp_1132_1 <= 0;
    end else begin
      if(_myaxi_write_req_fifo_enq && !_myaxi_write_req_fifo_full && (_myaxi_write_req_fifo_deq && !_myaxi_write_req_fifo_empty)) begin
        count__myaxi_write_req_fifo <= count__myaxi_write_req_fifo;
      end else if(_myaxi_write_req_fifo_enq && !_myaxi_write_req_fifo_full) begin
        count__myaxi_write_req_fifo <= count__myaxi_write_req_fifo + 1;
      end else if(_myaxi_write_req_fifo_deq && !_myaxi_write_req_fifo_empty) begin
        count__myaxi_write_req_fifo <= count__myaxi_write_req_fifo - 1;
      end 
      __tmp_1112_1 <= _tmp_1112;
      __tmp_1132_1 <= _tmp_1132;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_187_1 <= 0;
    end else begin
      __tmp_187_1 <= _tmp_187;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_190_1 <= 0;
    end else begin
      __tmp_190_1 <= _tmp_190;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_193_1 <= 0;
    end else begin
      __tmp_193_1 <= _tmp_193;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_196_1 <= 0;
    end else begin
      __tmp_196_1 <= _tmp_196;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_199_1 <= 0;
    end else begin
      __tmp_199_1 <= _tmp_199;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_202_1 <= 0;
    end else begin
      __tmp_202_1 <= _tmp_202;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_205_1 <= 0;
    end else begin
      __tmp_205_1 <= _tmp_205;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_208_1 <= 0;
    end else begin
      __tmp_208_1 <= _tmp_208;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_211_1 <= 0;
    end else begin
      __tmp_211_1 <= _tmp_211;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_214_1 <= 0;
    end else begin
      __tmp_214_1 <= _tmp_214;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_217_1 <= 0;
    end else begin
      __tmp_217_1 <= _tmp_217;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_220_1 <= 0;
    end else begin
      __tmp_220_1 <= _tmp_220;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_223_1 <= 0;
    end else begin
      __tmp_223_1 <= _tmp_223;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_226_1 <= 0;
    end else begin
      __tmp_226_1 <= _tmp_226;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_229_1 <= 0;
    end else begin
      __tmp_229_1 <= _tmp_229;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_232_1 <= 0;
    end else begin
      __tmp_232_1 <= _tmp_232;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_235_1 <= 0;
    end else begin
      __tmp_235_1 <= _tmp_235;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_238_1 <= 0;
    end else begin
      __tmp_238_1 <= _tmp_238;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_241_1 <= 0;
    end else begin
      __tmp_241_1 <= _tmp_241;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_244_1 <= 0;
    end else begin
      __tmp_244_1 <= _tmp_244;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_247_1 <= 0;
    end else begin
      __tmp_247_1 <= _tmp_247;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_250_1 <= 0;
    end else begin
      __tmp_250_1 <= _tmp_250;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_253_1 <= 0;
    end else begin
      __tmp_253_1 <= _tmp_253;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_256_1 <= 0;
    end else begin
      __tmp_256_1 <= _tmp_256;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_259_1 <= 0;
    end else begin
      __tmp_259_1 <= _tmp_259;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_262_1 <= 0;
    end else begin
      __tmp_262_1 <= _tmp_262;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_265_1 <= 0;
    end else begin
      __tmp_265_1 <= _tmp_265;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_268_1 <= 0;
    end else begin
      __tmp_268_1 <= _tmp_268;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_271_1 <= 0;
    end else begin
      __tmp_271_1 <= _tmp_271;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_274_1 <= 0;
    end else begin
      __tmp_274_1 <= _tmp_274;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_277_1 <= 0;
    end else begin
      __tmp_277_1 <= _tmp_277;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_280_1 <= 0;
    end else begin
      __tmp_280_1 <= _tmp_280;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_283_1 <= 0;
    end else begin
      __tmp_283_1 <= _tmp_283;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_286_1 <= 0;
    end else begin
      __tmp_286_1 <= _tmp_286;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_289_1 <= 0;
    end else begin
      __tmp_289_1 <= _tmp_289;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_292_1 <= 0;
    end else begin
      __tmp_292_1 <= _tmp_292;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_295_1 <= 0;
    end else begin
      __tmp_295_1 <= _tmp_295;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_298_1 <= 0;
    end else begin
      __tmp_298_1 <= _tmp_298;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_301_1 <= 0;
    end else begin
      __tmp_301_1 <= _tmp_301;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_304_1 <= 0;
    end else begin
      __tmp_304_1 <= _tmp_304;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_307_1 <= 0;
    end else begin
      __tmp_307_1 <= _tmp_307;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_310_1 <= 0;
    end else begin
      __tmp_310_1 <= _tmp_310;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_313_1 <= 0;
    end else begin
      __tmp_313_1 <= _tmp_313;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_316_1 <= 0;
    end else begin
      __tmp_316_1 <= _tmp_316;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_319_1 <= 0;
    end else begin
      __tmp_319_1 <= _tmp_319;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_322_1 <= 0;
    end else begin
      __tmp_322_1 <= _tmp_322;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_325_1 <= 0;
    end else begin
      __tmp_325_1 <= _tmp_325;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_328_1 <= 0;
    end else begin
      __tmp_328_1 <= _tmp_328;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_331_1 <= 0;
    end else begin
      __tmp_331_1 <= _tmp_331;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_334_1 <= 0;
    end else begin
      __tmp_334_1 <= _tmp_334;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_337_1 <= 0;
    end else begin
      __tmp_337_1 <= _tmp_337;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_340_1 <= 0;
    end else begin
      __tmp_340_1 <= _tmp_340;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_343_1 <= 0;
    end else begin
      __tmp_343_1 <= _tmp_343;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_346_1 <= 0;
    end else begin
      __tmp_346_1 <= _tmp_346;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_349_1 <= 0;
    end else begin
      __tmp_349_1 <= _tmp_349;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_352_1 <= 0;
    end else begin
      __tmp_352_1 <= _tmp_352;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_355_1 <= 0;
    end else begin
      __tmp_355_1 <= _tmp_355;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_358_1 <= 0;
    end else begin
      __tmp_358_1 <= _tmp_358;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_361_1 <= 0;
    end else begin
      __tmp_361_1 <= _tmp_361;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_364_1 <= 0;
    end else begin
      __tmp_364_1 <= _tmp_364;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_367_1 <= 0;
    end else begin
      __tmp_367_1 <= _tmp_367;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_370_1 <= 0;
    end else begin
      __tmp_370_1 <= _tmp_370;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_373_1 <= 0;
    end else begin
      __tmp_373_1 <= _tmp_373;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_376_1 <= 0;
    end else begin
      __tmp_376_1 <= _tmp_376;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1220_1 <= 0;
      __tmp_1289_1 <= 0;
    end else begin
      __tmp_1220_1 <= _tmp_1220;
      __tmp_1289_1 <= _tmp_1289;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1222_1 <= 0;
      __tmp_1291_1 <= 0;
    end else begin
      __tmp_1222_1 <= _tmp_1222;
      __tmp_1291_1 <= _tmp_1291;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1224_1 <= 0;
      __tmp_1293_1 <= 0;
    end else begin
      __tmp_1224_1 <= _tmp_1224;
      __tmp_1293_1 <= _tmp_1293;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1226_1 <= 0;
      __tmp_1295_1 <= 0;
    end else begin
      __tmp_1226_1 <= _tmp_1226;
      __tmp_1295_1 <= _tmp_1295;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1228_1 <= 0;
      __tmp_1297_1 <= 0;
    end else begin
      __tmp_1228_1 <= _tmp_1228;
      __tmp_1297_1 <= _tmp_1297;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1230_1 <= 0;
      __tmp_1299_1 <= 0;
    end else begin
      __tmp_1230_1 <= _tmp_1230;
      __tmp_1299_1 <= _tmp_1299;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1232_1 <= 0;
      __tmp_1301_1 <= 0;
    end else begin
      __tmp_1232_1 <= _tmp_1232;
      __tmp_1301_1 <= _tmp_1301;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1234_1 <= 0;
      __tmp_1303_1 <= 0;
    end else begin
      __tmp_1234_1 <= _tmp_1234;
      __tmp_1303_1 <= _tmp_1303;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1236_1 <= 0;
      __tmp_1305_1 <= 0;
    end else begin
      __tmp_1236_1 <= _tmp_1236;
      __tmp_1305_1 <= _tmp_1305;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1238_1 <= 0;
      __tmp_1307_1 <= 0;
    end else begin
      __tmp_1238_1 <= _tmp_1238;
      __tmp_1307_1 <= _tmp_1307;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1240_1 <= 0;
      __tmp_1309_1 <= 0;
    end else begin
      __tmp_1240_1 <= _tmp_1240;
      __tmp_1309_1 <= _tmp_1309;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1242_1 <= 0;
      __tmp_1311_1 <= 0;
    end else begin
      __tmp_1242_1 <= _tmp_1242;
      __tmp_1311_1 <= _tmp_1311;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1244_1 <= 0;
      __tmp_1313_1 <= 0;
    end else begin
      __tmp_1244_1 <= _tmp_1244;
      __tmp_1313_1 <= _tmp_1313;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1246_1 <= 0;
      __tmp_1315_1 <= 0;
    end else begin
      __tmp_1246_1 <= _tmp_1246;
      __tmp_1315_1 <= _tmp_1315;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1248_1 <= 0;
      __tmp_1317_1 <= 0;
    end else begin
      __tmp_1248_1 <= _tmp_1248;
      __tmp_1317_1 <= _tmp_1317;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1250_1 <= 0;
      __tmp_1319_1 <= 0;
    end else begin
      __tmp_1250_1 <= _tmp_1250;
      __tmp_1319_1 <= _tmp_1319;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1252_1 <= 0;
      __tmp_1321_1 <= 0;
    end else begin
      __tmp_1252_1 <= _tmp_1252;
      __tmp_1321_1 <= _tmp_1321;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1254_1 <= 0;
      __tmp_1323_1 <= 0;
    end else begin
      __tmp_1254_1 <= _tmp_1254;
      __tmp_1323_1 <= _tmp_1323;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1256_1 <= 0;
      __tmp_1325_1 <= 0;
    end else begin
      __tmp_1256_1 <= _tmp_1256;
      __tmp_1325_1 <= _tmp_1325;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1258_1 <= 0;
      __tmp_1327_1 <= 0;
    end else begin
      __tmp_1258_1 <= _tmp_1258;
      __tmp_1327_1 <= _tmp_1327;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1260_1 <= 0;
      __tmp_1329_1 <= 0;
    end else begin
      __tmp_1260_1 <= _tmp_1260;
      __tmp_1329_1 <= _tmp_1329;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1262_1 <= 0;
      __tmp_1331_1 <= 0;
    end else begin
      __tmp_1262_1 <= _tmp_1262;
      __tmp_1331_1 <= _tmp_1331;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1264_1 <= 0;
      __tmp_1333_1 <= 0;
    end else begin
      __tmp_1264_1 <= _tmp_1264;
      __tmp_1333_1 <= _tmp_1333;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1266_1 <= 0;
      __tmp_1335_1 <= 0;
    end else begin
      __tmp_1266_1 <= _tmp_1266;
      __tmp_1335_1 <= _tmp_1335;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1268_1 <= 0;
      __tmp_1337_1 <= 0;
    end else begin
      __tmp_1268_1 <= _tmp_1268;
      __tmp_1337_1 <= _tmp_1337;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1270_1 <= 0;
      __tmp_1339_1 <= 0;
    end else begin
      __tmp_1270_1 <= _tmp_1270;
      __tmp_1339_1 <= _tmp_1339;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1272_1 <= 0;
      __tmp_1341_1 <= 0;
    end else begin
      __tmp_1272_1 <= _tmp_1272;
      __tmp_1341_1 <= _tmp_1341;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1274_1 <= 0;
      __tmp_1343_1 <= 0;
    end else begin
      __tmp_1274_1 <= _tmp_1274;
      __tmp_1343_1 <= _tmp_1343;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1276_1 <= 0;
      __tmp_1345_1 <= 0;
    end else begin
      __tmp_1276_1 <= _tmp_1276;
      __tmp_1345_1 <= _tmp_1345;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1278_1 <= 0;
      __tmp_1347_1 <= 0;
    end else begin
      __tmp_1278_1 <= _tmp_1278;
      __tmp_1347_1 <= _tmp_1347;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1280_1 <= 0;
      __tmp_1349_1 <= 0;
    end else begin
      __tmp_1280_1 <= _tmp_1280;
      __tmp_1349_1 <= _tmp_1349;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1282_1 <= 0;
      __tmp_1351_1 <= 0;
    end else begin
      __tmp_1282_1 <= _tmp_1282;
      __tmp_1351_1 <= _tmp_1351;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1098_1 <= 0;
    end else begin
      __tmp_1098_1 <= _tmp_1098;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1101_1 <= 0;
    end else begin
      __tmp_1101_1 <= _tmp_1101;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      __tmp_1139_1 <= 0;
    end else begin
      __tmp_1139_1 <= _tmp_1139;
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _mystream_a0_source_ram_renable <= 0;
      _mystream_a0_source_fifo_deq <= 0;
      _mystream_a0_idle <= 1;
      _mystream_a1_source_ram_renable <= 0;
      _mystream_a1_source_fifo_deq <= 0;
      _mystream_a1_idle <= 1;
      _mystream_a2_source_ram_renable <= 0;
      _mystream_a2_source_fifo_deq <= 0;
      _mystream_a2_idle <= 1;
      _mystream_a3_source_ram_renable <= 0;
      _mystream_a3_source_fifo_deq <= 0;
      _mystream_a3_idle <= 1;
      _mystream_a4_source_ram_renable <= 0;
      _mystream_a4_source_fifo_deq <= 0;
      _mystream_a4_idle <= 1;
      _mystream_a5_source_ram_renable <= 0;
      _mystream_a5_source_fifo_deq <= 0;
      _mystream_a5_idle <= 1;
      _mystream_a6_source_ram_renable <= 0;
      _mystream_a6_source_fifo_deq <= 0;
      _mystream_a6_idle <= 1;
      _mystream_a7_source_ram_renable <= 0;
      _mystream_a7_source_fifo_deq <= 0;
      _mystream_a7_idle <= 1;
      _mystream_a8_source_ram_renable <= 0;
      _mystream_a8_source_fifo_deq <= 0;
      _mystream_a8_idle <= 1;
      _mystream_a9_source_ram_renable <= 0;
      _mystream_a9_source_fifo_deq <= 0;
      _mystream_a9_idle <= 1;
      _mystream_a10_source_ram_renable <= 0;
      _mystream_a10_source_fifo_deq <= 0;
      _mystream_a10_idle <= 1;
      _mystream_a11_source_ram_renable <= 0;
      _mystream_a11_source_fifo_deq <= 0;
      _mystream_a11_idle <= 1;
      _mystream_a12_source_ram_renable <= 0;
      _mystream_a12_source_fifo_deq <= 0;
      _mystream_a12_idle <= 1;
      _mystream_a13_source_ram_renable <= 0;
      _mystream_a13_source_fifo_deq <= 0;
      _mystream_a13_idle <= 1;
      _mystream_a14_source_ram_renable <= 0;
      _mystream_a14_source_fifo_deq <= 0;
      _mystream_a14_idle <= 1;
      _mystream_a15_source_ram_renable <= 0;
      _mystream_a15_source_fifo_deq <= 0;
      _mystream_a15_idle <= 1;
      _mystream_a16_source_ram_renable <= 0;
      _mystream_a16_source_fifo_deq <= 0;
      _mystream_a16_idle <= 1;
      _mystream_a17_source_ram_renable <= 0;
      _mystream_a17_source_fifo_deq <= 0;
      _mystream_a17_idle <= 1;
      _mystream_a18_source_ram_renable <= 0;
      _mystream_a18_source_fifo_deq <= 0;
      _mystream_a18_idle <= 1;
      _mystream_a19_source_ram_renable <= 0;
      _mystream_a19_source_fifo_deq <= 0;
      _mystream_a19_idle <= 1;
      _mystream_a20_source_ram_renable <= 0;
      _mystream_a20_source_fifo_deq <= 0;
      _mystream_a20_idle <= 1;
      _mystream_a21_source_ram_renable <= 0;
      _mystream_a21_source_fifo_deq <= 0;
      _mystream_a21_idle <= 1;
      _mystream_a22_source_ram_renable <= 0;
      _mystream_a22_source_fifo_deq <= 0;
      _mystream_a22_idle <= 1;
      _mystream_a23_source_ram_renable <= 0;
      _mystream_a23_source_fifo_deq <= 0;
      _mystream_a23_idle <= 1;
      _mystream_a24_source_ram_renable <= 0;
      _mystream_a24_source_fifo_deq <= 0;
      _mystream_a24_idle <= 1;
      _mystream_a25_source_ram_renable <= 0;
      _mystream_a25_source_fifo_deq <= 0;
      _mystream_a25_idle <= 1;
      _mystream_a26_source_ram_renable <= 0;
      _mystream_a26_source_fifo_deq <= 0;
      _mystream_a26_idle <= 1;
      _mystream_a27_source_ram_renable <= 0;
      _mystream_a27_source_fifo_deq <= 0;
      _mystream_a27_idle <= 1;
      _mystream_a28_source_ram_renable <= 0;
      _mystream_a28_source_fifo_deq <= 0;
      _mystream_a28_idle <= 1;
      _mystream_a29_source_ram_renable <= 0;
      _mystream_a29_source_fifo_deq <= 0;
      _mystream_a29_idle <= 1;
      _mystream_a30_source_ram_renable <= 0;
      _mystream_a30_source_fifo_deq <= 0;
      _mystream_a30_idle <= 1;
      _mystream_a31_source_ram_renable <= 0;
      _mystream_a31_source_fifo_deq <= 0;
      _mystream_a31_idle <= 1;
      _mystream_b0_source_ram_renable <= 0;
      _mystream_b0_source_fifo_deq <= 0;
      _mystream_b0_idle <= 1;
      _mystream_b1_source_ram_renable <= 0;
      _mystream_b1_source_fifo_deq <= 0;
      _mystream_b1_idle <= 1;
      _mystream_b2_source_ram_renable <= 0;
      _mystream_b2_source_fifo_deq <= 0;
      _mystream_b2_idle <= 1;
      _mystream_b3_source_ram_renable <= 0;
      _mystream_b3_source_fifo_deq <= 0;
      _mystream_b3_idle <= 1;
      _mystream_b4_source_ram_renable <= 0;
      _mystream_b4_source_fifo_deq <= 0;
      _mystream_b4_idle <= 1;
      _mystream_b5_source_ram_renable <= 0;
      _mystream_b5_source_fifo_deq <= 0;
      _mystream_b5_idle <= 1;
      _mystream_b6_source_ram_renable <= 0;
      _mystream_b6_source_fifo_deq <= 0;
      _mystream_b6_idle <= 1;
      _mystream_b7_source_ram_renable <= 0;
      _mystream_b7_source_fifo_deq <= 0;
      _mystream_b7_idle <= 1;
      _mystream_b8_source_ram_renable <= 0;
      _mystream_b8_source_fifo_deq <= 0;
      _mystream_b8_idle <= 1;
      _mystream_b9_source_ram_renable <= 0;
      _mystream_b9_source_fifo_deq <= 0;
      _mystream_b9_idle <= 1;
      _mystream_b10_source_ram_renable <= 0;
      _mystream_b10_source_fifo_deq <= 0;
      _mystream_b10_idle <= 1;
      _mystream_b11_source_ram_renable <= 0;
      _mystream_b11_source_fifo_deq <= 0;
      _mystream_b11_idle <= 1;
      _mystream_b12_source_ram_renable <= 0;
      _mystream_b12_source_fifo_deq <= 0;
      _mystream_b12_idle <= 1;
      _mystream_b13_source_ram_renable <= 0;
      _mystream_b13_source_fifo_deq <= 0;
      _mystream_b13_idle <= 1;
      _mystream_b14_source_ram_renable <= 0;
      _mystream_b14_source_fifo_deq <= 0;
      _mystream_b14_idle <= 1;
      _mystream_b15_source_ram_renable <= 0;
      _mystream_b15_source_fifo_deq <= 0;
      _mystream_b15_idle <= 1;
      _mystream_b16_source_ram_renable <= 0;
      _mystream_b16_source_fifo_deq <= 0;
      _mystream_b16_idle <= 1;
      _mystream_b17_source_ram_renable <= 0;
      _mystream_b17_source_fifo_deq <= 0;
      _mystream_b17_idle <= 1;
      _mystream_b18_source_ram_renable <= 0;
      _mystream_b18_source_fifo_deq <= 0;
      _mystream_b18_idle <= 1;
      _mystream_b19_source_ram_renable <= 0;
      _mystream_b19_source_fifo_deq <= 0;
      _mystream_b19_idle <= 1;
      _mystream_b20_source_ram_renable <= 0;
      _mystream_b20_source_fifo_deq <= 0;
      _mystream_b20_idle <= 1;
      _mystream_b21_source_ram_renable <= 0;
      _mystream_b21_source_fifo_deq <= 0;
      _mystream_b21_idle <= 1;
      _mystream_b22_source_ram_renable <= 0;
      _mystream_b22_source_fifo_deq <= 0;
      _mystream_b22_idle <= 1;
      _mystream_b23_source_ram_renable <= 0;
      _mystream_b23_source_fifo_deq <= 0;
      _mystream_b23_idle <= 1;
      _mystream_b24_source_ram_renable <= 0;
      _mystream_b24_source_fifo_deq <= 0;
      _mystream_b24_idle <= 1;
      _mystream_b25_source_ram_renable <= 0;
      _mystream_b25_source_fifo_deq <= 0;
      _mystream_b25_idle <= 1;
      _mystream_b26_source_ram_renable <= 0;
      _mystream_b26_source_fifo_deq <= 0;
      _mystream_b26_idle <= 1;
      _mystream_b27_source_ram_renable <= 0;
      _mystream_b27_source_fifo_deq <= 0;
      _mystream_b27_idle <= 1;
      _mystream_b28_source_ram_renable <= 0;
      _mystream_b28_source_fifo_deq <= 0;
      _mystream_b28_idle <= 1;
      _mystream_b29_source_ram_renable <= 0;
      _mystream_b29_source_fifo_deq <= 0;
      _mystream_b29_idle <= 1;
      _mystream_b30_source_ram_renable <= 0;
      _mystream_b30_source_fifo_deq <= 0;
      _mystream_b30_idle <= 1;
      _mystream_b31_source_ram_renable <= 0;
      _mystream_b31_source_fifo_deq <= 0;
      _mystream_b31_idle <= 1;
      _mystream_bias0_source_ram_renable <= 0;
      _mystream_bias0_source_fifo_deq <= 0;
      _mystream_bias0_idle <= 1;
      _mystream_bias1_source_ram_renable <= 0;
      _mystream_bias1_source_fifo_deq <= 0;
      _mystream_bias1_idle <= 1;
      _mystream_bias2_source_ram_renable <= 0;
      _mystream_bias2_source_fifo_deq <= 0;
      _mystream_bias2_idle <= 1;
      _mystream_bias3_source_ram_renable <= 0;
      _mystream_bias3_source_fifo_deq <= 0;
      _mystream_bias3_idle <= 1;
      _mystream_bias4_source_ram_renable <= 0;
      _mystream_bias4_source_fifo_deq <= 0;
      _mystream_bias4_idle <= 1;
      _mystream_bias5_source_ram_renable <= 0;
      _mystream_bias5_source_fifo_deq <= 0;
      _mystream_bias5_idle <= 1;
      _mystream_bias6_source_ram_renable <= 0;
      _mystream_bias6_source_fifo_deq <= 0;
      _mystream_bias6_idle <= 1;
      _mystream_bias7_source_ram_renable <= 0;
      _mystream_bias7_source_fifo_deq <= 0;
      _mystream_bias7_idle <= 1;
      _mystream_bias8_source_ram_renable <= 0;
      _mystream_bias8_source_fifo_deq <= 0;
      _mystream_bias8_idle <= 1;
      _mystream_bias9_source_ram_renable <= 0;
      _mystream_bias9_source_fifo_deq <= 0;
      _mystream_bias9_idle <= 1;
      _mystream_bias10_source_ram_renable <= 0;
      _mystream_bias10_source_fifo_deq <= 0;
      _mystream_bias10_idle <= 1;
      _mystream_bias11_source_ram_renable <= 0;
      _mystream_bias11_source_fifo_deq <= 0;
      _mystream_bias11_idle <= 1;
      _mystream_bias12_source_ram_renable <= 0;
      _mystream_bias12_source_fifo_deq <= 0;
      _mystream_bias12_idle <= 1;
      _mystream_bias13_source_ram_renable <= 0;
      _mystream_bias13_source_fifo_deq <= 0;
      _mystream_bias13_idle <= 1;
      _mystream_bias14_source_ram_renable <= 0;
      _mystream_bias14_source_fifo_deq <= 0;
      _mystream_bias14_idle <= 1;
      _mystream_bias15_source_ram_renable <= 0;
      _mystream_bias15_source_fifo_deq <= 0;
      _mystream_bias15_idle <= 1;
      _mystream_bias16_source_ram_renable <= 0;
      _mystream_bias16_source_fifo_deq <= 0;
      _mystream_bias16_idle <= 1;
      _mystream_bias17_source_ram_renable <= 0;
      _mystream_bias17_source_fifo_deq <= 0;
      _mystream_bias17_idle <= 1;
      _mystream_bias18_source_ram_renable <= 0;
      _mystream_bias18_source_fifo_deq <= 0;
      _mystream_bias18_idle <= 1;
      _mystream_bias19_source_ram_renable <= 0;
      _mystream_bias19_source_fifo_deq <= 0;
      _mystream_bias19_idle <= 1;
      _mystream_bias20_source_ram_renable <= 0;
      _mystream_bias20_source_fifo_deq <= 0;
      _mystream_bias20_idle <= 1;
      _mystream_bias21_source_ram_renable <= 0;
      _mystream_bias21_source_fifo_deq <= 0;
      _mystream_bias21_idle <= 1;
      _mystream_bias22_source_ram_renable <= 0;
      _mystream_bias22_source_fifo_deq <= 0;
      _mystream_bias22_idle <= 1;
      _mystream_bias23_source_ram_renable <= 0;
      _mystream_bias23_source_fifo_deq <= 0;
      _mystream_bias23_idle <= 1;
      _mystream_bias24_source_ram_renable <= 0;
      _mystream_bias24_source_fifo_deq <= 0;
      _mystream_bias24_idle <= 1;
      _mystream_bias25_source_ram_renable <= 0;
      _mystream_bias25_source_fifo_deq <= 0;
      _mystream_bias25_idle <= 1;
      _mystream_bias26_source_ram_renable <= 0;
      _mystream_bias26_source_fifo_deq <= 0;
      _mystream_bias26_idle <= 1;
      _mystream_bias27_source_ram_renable <= 0;
      _mystream_bias27_source_fifo_deq <= 0;
      _mystream_bias27_idle <= 1;
      _mystream_bias28_source_ram_renable <= 0;
      _mystream_bias28_source_fifo_deq <= 0;
      _mystream_bias28_idle <= 1;
      _mystream_bias29_source_ram_renable <= 0;
      _mystream_bias29_source_fifo_deq <= 0;
      _mystream_bias29_idle <= 1;
      _mystream_bias30_source_ram_renable <= 0;
      _mystream_bias30_source_fifo_deq <= 0;
      _mystream_bias30_idle <= 1;
      _mystream_bias31_source_ram_renable <= 0;
      _mystream_bias31_source_fifo_deq <= 0;
      _mystream_bias31_idle <= 1;
      _mystream_sum_vec0_sink_wenable <= 0;
      _mystream_sum_vec0_sink_fifo_enq <= 0;
      _mystream_sum_vec1_sink_wenable <= 0;
      _mystream_sum_vec1_sink_fifo_enq <= 0;
      _mystream_sum_vec2_sink_wenable <= 0;
      _mystream_sum_vec2_sink_fifo_enq <= 0;
      _mystream_sum_vec3_sink_wenable <= 0;
      _mystream_sum_vec3_sink_fifo_enq <= 0;
      _mystream_sum_vec4_sink_wenable <= 0;
      _mystream_sum_vec4_sink_fifo_enq <= 0;
      _mystream_sum_vec5_sink_wenable <= 0;
      _mystream_sum_vec5_sink_fifo_enq <= 0;
      _mystream_sum_vec6_sink_wenable <= 0;
      _mystream_sum_vec6_sink_fifo_enq <= 0;
      _mystream_sum_vec7_sink_wenable <= 0;
      _mystream_sum_vec7_sink_fifo_enq <= 0;
      _mystream_sum_vec8_sink_wenable <= 0;
      _mystream_sum_vec8_sink_fifo_enq <= 0;
      _mystream_sum_vec9_sink_wenable <= 0;
      _mystream_sum_vec9_sink_fifo_enq <= 0;
      _mystream_sum_vec10_sink_wenable <= 0;
      _mystream_sum_vec10_sink_fifo_enq <= 0;
      _mystream_sum_vec11_sink_wenable <= 0;
      _mystream_sum_vec11_sink_fifo_enq <= 0;
      _mystream_sum_vec12_sink_wenable <= 0;
      _mystream_sum_vec12_sink_fifo_enq <= 0;
      _mystream_sum_vec13_sink_wenable <= 0;
      _mystream_sum_vec13_sink_fifo_enq <= 0;
      _mystream_sum_vec14_sink_wenable <= 0;
      _mystream_sum_vec14_sink_fifo_enq <= 0;
      _mystream_sum_vec15_sink_wenable <= 0;
      _mystream_sum_vec15_sink_fifo_enq <= 0;
      _mystream_sum_vec16_sink_wenable <= 0;
      _mystream_sum_vec16_sink_fifo_enq <= 0;
      _mystream_sum_vec17_sink_wenable <= 0;
      _mystream_sum_vec17_sink_fifo_enq <= 0;
      _mystream_sum_vec18_sink_wenable <= 0;
      _mystream_sum_vec18_sink_fifo_enq <= 0;
      _mystream_sum_vec19_sink_wenable <= 0;
      _mystream_sum_vec19_sink_fifo_enq <= 0;
      _mystream_sum_vec20_sink_wenable <= 0;
      _mystream_sum_vec20_sink_fifo_enq <= 0;
      _mystream_sum_vec21_sink_wenable <= 0;
      _mystream_sum_vec21_sink_fifo_enq <= 0;
      _mystream_sum_vec22_sink_wenable <= 0;
      _mystream_sum_vec22_sink_fifo_enq <= 0;
      _mystream_sum_vec23_sink_wenable <= 0;
      _mystream_sum_vec23_sink_fifo_enq <= 0;
      _mystream_sum_vec24_sink_wenable <= 0;
      _mystream_sum_vec24_sink_fifo_enq <= 0;
      _mystream_sum_vec25_sink_wenable <= 0;
      _mystream_sum_vec25_sink_fifo_enq <= 0;
      _mystream_sum_vec26_sink_wenable <= 0;
      _mystream_sum_vec26_sink_fifo_enq <= 0;
      _mystream_sum_vec27_sink_wenable <= 0;
      _mystream_sum_vec27_sink_fifo_enq <= 0;
      _mystream_sum_vec28_sink_wenable <= 0;
      _mystream_sum_vec28_sink_fifo_enq <= 0;
      _mystream_sum_vec29_sink_wenable <= 0;
      _mystream_sum_vec29_sink_fifo_enq <= 0;
      _mystream_sum_vec30_sink_wenable <= 0;
      _mystream_sum_vec30_sink_fifo_enq <= 0;
      _mystream_sum_vec31_sink_wenable <= 0;
      _mystream_sum_vec31_sink_fifo_enq <= 0;
      __mystream_stream_ivalid_1 <= 0;
      __mystream_stream_ivalid_2 <= 0;
      __mystream_stream_ivalid_3 <= 0;
      __mystream_stream_ivalid_4 <= 0;
      _plus_data_98 <= 0;
      _plus_data_99 <= 0;
      _plus_data_100 <= 0;
      _plus_data_101 <= 0;
      _plus_data_102 <= 0;
      _plus_data_103 <= 0;
      _plus_data_104 <= 0;
      _plus_data_105 <= 0;
      _plus_data_106 <= 0;
      _plus_data_107 <= 0;
      _plus_data_108 <= 0;
      _plus_data_109 <= 0;
      _plus_data_110 <= 0;
      _plus_data_111 <= 0;
      _plus_data_112 <= 0;
      _plus_data_113 <= 0;
      _plus_data_114 <= 0;
      _plus_data_115 <= 0;
      _plus_data_116 <= 0;
      _plus_data_117 <= 0;
      _plus_data_118 <= 0;
      _plus_data_119 <= 0;
      _plus_data_120 <= 0;
      _plus_data_121 <= 0;
      _plus_data_122 <= 0;
      _plus_data_123 <= 0;
      _plus_data_124 <= 0;
      _plus_data_125 <= 0;
      _plus_data_126 <= 0;
      _plus_data_127 <= 0;
      _plus_data_128 <= 0;
      _plus_data_129 <= 0;
      _counter_data_131 <= 1'sd0;
      _counter_count_131 <= 1'sd0;
      __delay_data_294__variable_1 <= 0;
      _plus_data_134 <= 0;
      _plus_data_137 <= 0;
      _plus_data_140 <= 0;
      _plus_data_143 <= 0;
      _plus_data_146 <= 0;
      _plus_data_149 <= 0;
      _plus_data_152 <= 0;
      _plus_data_155 <= 0;
      _plus_data_158 <= 0;
      _plus_data_161 <= 0;
      _plus_data_164 <= 0;
      _plus_data_167 <= 0;
      _plus_data_170 <= 0;
      _plus_data_173 <= 0;
      _plus_data_176 <= 0;
      _plus_data_179 <= 0;
      _plus_data_182 <= 0;
      _plus_data_185 <= 0;
      _plus_data_188 <= 0;
      _plus_data_191 <= 0;
      _plus_data_194 <= 0;
      _plus_data_197 <= 0;
      _plus_data_200 <= 0;
      _plus_data_203 <= 0;
      _plus_data_206 <= 0;
      _plus_data_209 <= 0;
      _plus_data_212 <= 0;
      _plus_data_215 <= 0;
      _plus_data_218 <= 0;
      _plus_data_221 <= 0;
      _plus_data_224 <= 0;
      _plus_data_227 <= 0;
      __delay_data_295__delay_294__variable_1 <= 0;
      __delay_data_296_plus_98 <= 0;
      __delay_data_298_plus_99 <= 0;
      __delay_data_300_plus_100 <= 0;
      __delay_data_302_plus_101 <= 0;
      __delay_data_304_plus_102 <= 0;
      __delay_data_306_plus_103 <= 0;
      __delay_data_308_plus_104 <= 0;
      __delay_data_310_plus_105 <= 0;
      __delay_data_312_plus_106 <= 0;
      __delay_data_314_plus_107 <= 0;
      __delay_data_316_plus_108 <= 0;
      __delay_data_318_plus_109 <= 0;
      __delay_data_320_plus_110 <= 0;
      __delay_data_322_plus_111 <= 0;
      __delay_data_324_plus_112 <= 0;
      __delay_data_326_plus_113 <= 0;
      __delay_data_328_plus_114 <= 0;
      __delay_data_330_plus_115 <= 0;
      __delay_data_332_plus_116 <= 0;
      __delay_data_334_plus_117 <= 0;
      __delay_data_336_plus_118 <= 0;
      __delay_data_338_plus_119 <= 0;
      __delay_data_340_plus_120 <= 0;
      __delay_data_342_plus_121 <= 0;
      __delay_data_344_plus_122 <= 0;
      __delay_data_346_plus_123 <= 0;
      __delay_data_348_plus_124 <= 0;
      __delay_data_350_plus_125 <= 0;
      __delay_data_352_plus_126 <= 0;
      __delay_data_354_plus_127 <= 0;
      __delay_data_356_plus_128 <= 0;
      __delay_data_358_plus_129 <= 0;
      _greatereq_data_136 <= 0;
      _greatereq_data_139 <= 0;
      _greatereq_data_142 <= 0;
      _greatereq_data_145 <= 0;
      _greatereq_data_148 <= 0;
      _greatereq_data_151 <= 0;
      _greatereq_data_154 <= 0;
      _greatereq_data_157 <= 0;
      _greatereq_data_160 <= 0;
      _greatereq_data_163 <= 0;
      _greatereq_data_166 <= 0;
      _greatereq_data_169 <= 0;
      _greatereq_data_172 <= 0;
      _greatereq_data_175 <= 0;
      _greatereq_data_178 <= 0;
      _greatereq_data_181 <= 0;
      _greatereq_data_184 <= 0;
      _greatereq_data_187 <= 0;
      _greatereq_data_190 <= 0;
      _greatereq_data_193 <= 0;
      _greatereq_data_196 <= 0;
      _greatereq_data_199 <= 0;
      _greatereq_data_202 <= 0;
      _greatereq_data_205 <= 0;
      _greatereq_data_208 <= 0;
      _greatereq_data_211 <= 0;
      _greatereq_data_214 <= 0;
      _greatereq_data_217 <= 0;
      _greatereq_data_220 <= 0;
      _greatereq_data_223 <= 0;
      _greatereq_data_226 <= 0;
      _greatereq_data_229 <= 0;
      __delay_data_297__delay_296_plus_98 <= 0;
      __delay_data_299__delay_298_plus_99 <= 0;
      __delay_data_301__delay_300_plus_100 <= 0;
      __delay_data_303__delay_302_plus_101 <= 0;
      __delay_data_305__delay_304_plus_102 <= 0;
      __delay_data_307__delay_306_plus_103 <= 0;
      __delay_data_309__delay_308_plus_104 <= 0;
      __delay_data_311__delay_310_plus_105 <= 0;
      __delay_data_313__delay_312_plus_106 <= 0;
      __delay_data_315__delay_314_plus_107 <= 0;
      __delay_data_317__delay_316_plus_108 <= 0;
      __delay_data_319__delay_318_plus_109 <= 0;
      __delay_data_321__delay_320_plus_110 <= 0;
      __delay_data_323__delay_322_plus_111 <= 0;
      __delay_data_325__delay_324_plus_112 <= 0;
      __delay_data_327__delay_326_plus_113 <= 0;
      __delay_data_329__delay_328_plus_114 <= 0;
      __delay_data_331__delay_330_plus_115 <= 0;
      __delay_data_333__delay_332_plus_116 <= 0;
      __delay_data_335__delay_334_plus_117 <= 0;
      __delay_data_337__delay_336_plus_118 <= 0;
      __delay_data_339__delay_338_plus_119 <= 0;
      __delay_data_341__delay_340_plus_120 <= 0;
      __delay_data_343__delay_342_plus_121 <= 0;
      __delay_data_345__delay_344_plus_122 <= 0;
      __delay_data_347__delay_346_plus_123 <= 0;
      __delay_data_349__delay_348_plus_124 <= 0;
      __delay_data_351__delay_350_plus_125 <= 0;
      __delay_data_353__delay_352_plus_126 <= 0;
      __delay_data_355__delay_354_plus_127 <= 0;
      __delay_data_357__delay_356_plus_128 <= 0;
      __delay_data_359__delay_358_plus_129 <= 0;
      _cond_data_230 <= 0;
      _cond_data_232 <= 0;
      _cond_data_234 <= 0;
      _cond_data_236 <= 0;
      _cond_data_238 <= 0;
      _cond_data_240 <= 0;
      _cond_data_242 <= 0;
      _cond_data_244 <= 0;
      _cond_data_246 <= 0;
      _cond_data_248 <= 0;
      _cond_data_250 <= 0;
      _cond_data_252 <= 0;
      _cond_data_254 <= 0;
      _cond_data_256 <= 0;
      _cond_data_258 <= 0;
      _cond_data_260 <= 0;
      _cond_data_262 <= 0;
      _cond_data_264 <= 0;
      _cond_data_266 <= 0;
      _cond_data_268 <= 0;
      _cond_data_270 <= 0;
      _cond_data_272 <= 0;
      _cond_data_274 <= 0;
      _cond_data_276 <= 0;
      _cond_data_278 <= 0;
      _cond_data_280 <= 0;
      _cond_data_282 <= 0;
      _cond_data_284 <= 0;
      _cond_data_286 <= 0;
      _cond_data_288 <= 0;
      _cond_data_290 <= 0;
      _cond_data_292 <= 0;
      _mystream_tensor_size_next_parameter_data <= 0;
      __variable_wdata_1 <= 0;
      _mystream_size_next_parameter_data <= 0;
      __variable_wdata_0 <= 0;
      _mystream_a0_source_mode <= 5'b0;
      _mystream_a0_source_offset <= 0;
      _mystream_a0_source_size <= 0;
      _mystream_a0_source_stride <= 0;
      _mystream_a0_source_sel <= 0;
      _mystream_a0_source_offset_buf <= 0;
      _mystream_a0_source_size_buf <= 0;
      _mystream_a0_source_stride_buf <= 0;
      __variable_wdata_2 <= 0;
      _mystream_a0_source_ram_raddr <= 0;
      _mystream_a0_source_count <= 0;
      _mystream_a1_source_mode <= 5'b0;
      _mystream_a1_source_offset <= 0;
      _mystream_a1_source_size <= 0;
      _mystream_a1_source_stride <= 0;
      _mystream_a1_source_sel <= 0;
      _mystream_a1_source_offset_buf <= 0;
      _mystream_a1_source_size_buf <= 0;
      _mystream_a1_source_stride_buf <= 0;
      __variable_wdata_3 <= 0;
      _mystream_a1_source_ram_raddr <= 0;
      _mystream_a1_source_count <= 0;
      _mystream_a2_source_mode <= 5'b0;
      _mystream_a2_source_offset <= 0;
      _mystream_a2_source_size <= 0;
      _mystream_a2_source_stride <= 0;
      _mystream_a2_source_sel <= 0;
      _mystream_a2_source_offset_buf <= 0;
      _mystream_a2_source_size_buf <= 0;
      _mystream_a2_source_stride_buf <= 0;
      __variable_wdata_4 <= 0;
      _mystream_a2_source_ram_raddr <= 0;
      _mystream_a2_source_count <= 0;
      _mystream_a3_source_mode <= 5'b0;
      _mystream_a3_source_offset <= 0;
      _mystream_a3_source_size <= 0;
      _mystream_a3_source_stride <= 0;
      _mystream_a3_source_sel <= 0;
      _mystream_a3_source_offset_buf <= 0;
      _mystream_a3_source_size_buf <= 0;
      _mystream_a3_source_stride_buf <= 0;
      __variable_wdata_5 <= 0;
      _mystream_a3_source_ram_raddr <= 0;
      _mystream_a3_source_count <= 0;
      _mystream_a4_source_mode <= 5'b0;
      _mystream_a4_source_offset <= 0;
      _mystream_a4_source_size <= 0;
      _mystream_a4_source_stride <= 0;
      _mystream_a4_source_sel <= 0;
      _mystream_a4_source_offset_buf <= 0;
      _mystream_a4_source_size_buf <= 0;
      _mystream_a4_source_stride_buf <= 0;
      __variable_wdata_6 <= 0;
      _mystream_a4_source_ram_raddr <= 0;
      _mystream_a4_source_count <= 0;
      _mystream_a5_source_mode <= 5'b0;
      _mystream_a5_source_offset <= 0;
      _mystream_a5_source_size <= 0;
      _mystream_a5_source_stride <= 0;
      _mystream_a5_source_sel <= 0;
      _mystream_a5_source_offset_buf <= 0;
      _mystream_a5_source_size_buf <= 0;
      _mystream_a5_source_stride_buf <= 0;
      __variable_wdata_7 <= 0;
      _mystream_a5_source_ram_raddr <= 0;
      _mystream_a5_source_count <= 0;
      _mystream_a6_source_mode <= 5'b0;
      _mystream_a6_source_offset <= 0;
      _mystream_a6_source_size <= 0;
      _mystream_a6_source_stride <= 0;
      _mystream_a6_source_sel <= 0;
      _mystream_a6_source_offset_buf <= 0;
      _mystream_a6_source_size_buf <= 0;
      _mystream_a6_source_stride_buf <= 0;
      __variable_wdata_8 <= 0;
      _mystream_a6_source_ram_raddr <= 0;
      _mystream_a6_source_count <= 0;
      _mystream_a7_source_mode <= 5'b0;
      _mystream_a7_source_offset <= 0;
      _mystream_a7_source_size <= 0;
      _mystream_a7_source_stride <= 0;
      _mystream_a7_source_sel <= 0;
      _mystream_a7_source_offset_buf <= 0;
      _mystream_a7_source_size_buf <= 0;
      _mystream_a7_source_stride_buf <= 0;
      __variable_wdata_9 <= 0;
      _mystream_a7_source_ram_raddr <= 0;
      _mystream_a7_source_count <= 0;
      _mystream_a8_source_mode <= 5'b0;
      _mystream_a8_source_offset <= 0;
      _mystream_a8_source_size <= 0;
      _mystream_a8_source_stride <= 0;
      _mystream_a8_source_sel <= 0;
      _mystream_a8_source_offset_buf <= 0;
      _mystream_a8_source_size_buf <= 0;
      _mystream_a8_source_stride_buf <= 0;
      __variable_wdata_10 <= 0;
      _mystream_a8_source_ram_raddr <= 0;
      _mystream_a8_source_count <= 0;
      _mystream_a9_source_mode <= 5'b0;
      _mystream_a9_source_offset <= 0;
      _mystream_a9_source_size <= 0;
      _mystream_a9_source_stride <= 0;
      _mystream_a9_source_sel <= 0;
      _mystream_a9_source_offset_buf <= 0;
      _mystream_a9_source_size_buf <= 0;
      _mystream_a9_source_stride_buf <= 0;
      __variable_wdata_11 <= 0;
      _mystream_a9_source_ram_raddr <= 0;
      _mystream_a9_source_count <= 0;
      _mystream_a10_source_mode <= 5'b0;
      _mystream_a10_source_offset <= 0;
      _mystream_a10_source_size <= 0;
      _mystream_a10_source_stride <= 0;
      _mystream_a10_source_sel <= 0;
      _mystream_a10_source_offset_buf <= 0;
      _mystream_a10_source_size_buf <= 0;
      _mystream_a10_source_stride_buf <= 0;
      __variable_wdata_12 <= 0;
      _mystream_a10_source_ram_raddr <= 0;
      _mystream_a10_source_count <= 0;
      _mystream_a11_source_mode <= 5'b0;
      _mystream_a11_source_offset <= 0;
      _mystream_a11_source_size <= 0;
      _mystream_a11_source_stride <= 0;
      _mystream_a11_source_sel <= 0;
      _mystream_a11_source_offset_buf <= 0;
      _mystream_a11_source_size_buf <= 0;
      _mystream_a11_source_stride_buf <= 0;
      __variable_wdata_13 <= 0;
      _mystream_a11_source_ram_raddr <= 0;
      _mystream_a11_source_count <= 0;
      _mystream_a12_source_mode <= 5'b0;
      _mystream_a12_source_offset <= 0;
      _mystream_a12_source_size <= 0;
      _mystream_a12_source_stride <= 0;
      _mystream_a12_source_sel <= 0;
      _mystream_a12_source_offset_buf <= 0;
      _mystream_a12_source_size_buf <= 0;
      _mystream_a12_source_stride_buf <= 0;
      __variable_wdata_14 <= 0;
      _mystream_a12_source_ram_raddr <= 0;
      _mystream_a12_source_count <= 0;
      _mystream_a13_source_mode <= 5'b0;
      _mystream_a13_source_offset <= 0;
      _mystream_a13_source_size <= 0;
      _mystream_a13_source_stride <= 0;
      _mystream_a13_source_sel <= 0;
      _mystream_a13_source_offset_buf <= 0;
      _mystream_a13_source_size_buf <= 0;
      _mystream_a13_source_stride_buf <= 0;
      __variable_wdata_15 <= 0;
      _mystream_a13_source_ram_raddr <= 0;
      _mystream_a13_source_count <= 0;
      _mystream_a14_source_mode <= 5'b0;
      _mystream_a14_source_offset <= 0;
      _mystream_a14_source_size <= 0;
      _mystream_a14_source_stride <= 0;
      _mystream_a14_source_sel <= 0;
      _mystream_a14_source_offset_buf <= 0;
      _mystream_a14_source_size_buf <= 0;
      _mystream_a14_source_stride_buf <= 0;
      __variable_wdata_16 <= 0;
      _mystream_a14_source_ram_raddr <= 0;
      _mystream_a14_source_count <= 0;
      _mystream_a15_source_mode <= 5'b0;
      _mystream_a15_source_offset <= 0;
      _mystream_a15_source_size <= 0;
      _mystream_a15_source_stride <= 0;
      _mystream_a15_source_sel <= 0;
      _mystream_a15_source_offset_buf <= 0;
      _mystream_a15_source_size_buf <= 0;
      _mystream_a15_source_stride_buf <= 0;
      __variable_wdata_17 <= 0;
      _mystream_a15_source_ram_raddr <= 0;
      _mystream_a15_source_count <= 0;
      _mystream_a16_source_mode <= 5'b0;
      _mystream_a16_source_offset <= 0;
      _mystream_a16_source_size <= 0;
      _mystream_a16_source_stride <= 0;
      _mystream_a16_source_sel <= 0;
      _mystream_a16_source_offset_buf <= 0;
      _mystream_a16_source_size_buf <= 0;
      _mystream_a16_source_stride_buf <= 0;
      __variable_wdata_18 <= 0;
      _mystream_a16_source_ram_raddr <= 0;
      _mystream_a16_source_count <= 0;
      _mystream_a17_source_mode <= 5'b0;
      _mystream_a17_source_offset <= 0;
      _mystream_a17_source_size <= 0;
      _mystream_a17_source_stride <= 0;
      _mystream_a17_source_sel <= 0;
      _mystream_a17_source_offset_buf <= 0;
      _mystream_a17_source_size_buf <= 0;
      _mystream_a17_source_stride_buf <= 0;
      __variable_wdata_19 <= 0;
      _mystream_a17_source_ram_raddr <= 0;
      _mystream_a17_source_count <= 0;
      _mystream_a18_source_mode <= 5'b0;
      _mystream_a18_source_offset <= 0;
      _mystream_a18_source_size <= 0;
      _mystream_a18_source_stride <= 0;
      _mystream_a18_source_sel <= 0;
      _mystream_a18_source_offset_buf <= 0;
      _mystream_a18_source_size_buf <= 0;
      _mystream_a18_source_stride_buf <= 0;
      __variable_wdata_20 <= 0;
      _mystream_a18_source_ram_raddr <= 0;
      _mystream_a18_source_count <= 0;
      _mystream_a19_source_mode <= 5'b0;
      _mystream_a19_source_offset <= 0;
      _mystream_a19_source_size <= 0;
      _mystream_a19_source_stride <= 0;
      _mystream_a19_source_sel <= 0;
      _mystream_a19_source_offset_buf <= 0;
      _mystream_a19_source_size_buf <= 0;
      _mystream_a19_source_stride_buf <= 0;
      __variable_wdata_21 <= 0;
      _mystream_a19_source_ram_raddr <= 0;
      _mystream_a19_source_count <= 0;
      _mystream_a20_source_mode <= 5'b0;
      _mystream_a20_source_offset <= 0;
      _mystream_a20_source_size <= 0;
      _mystream_a20_source_stride <= 0;
      _mystream_a20_source_sel <= 0;
      _mystream_a20_source_offset_buf <= 0;
      _mystream_a20_source_size_buf <= 0;
      _mystream_a20_source_stride_buf <= 0;
      __variable_wdata_22 <= 0;
      _mystream_a20_source_ram_raddr <= 0;
      _mystream_a20_source_count <= 0;
      _mystream_a21_source_mode <= 5'b0;
      _mystream_a21_source_offset <= 0;
      _mystream_a21_source_size <= 0;
      _mystream_a21_source_stride <= 0;
      _mystream_a21_source_sel <= 0;
      _mystream_a21_source_offset_buf <= 0;
      _mystream_a21_source_size_buf <= 0;
      _mystream_a21_source_stride_buf <= 0;
      __variable_wdata_23 <= 0;
      _mystream_a21_source_ram_raddr <= 0;
      _mystream_a21_source_count <= 0;
      _mystream_a22_source_mode <= 5'b0;
      _mystream_a22_source_offset <= 0;
      _mystream_a22_source_size <= 0;
      _mystream_a22_source_stride <= 0;
      _mystream_a22_source_sel <= 0;
      _mystream_a22_source_offset_buf <= 0;
      _mystream_a22_source_size_buf <= 0;
      _mystream_a22_source_stride_buf <= 0;
      __variable_wdata_24 <= 0;
      _mystream_a22_source_ram_raddr <= 0;
      _mystream_a22_source_count <= 0;
      _mystream_a23_source_mode <= 5'b0;
      _mystream_a23_source_offset <= 0;
      _mystream_a23_source_size <= 0;
      _mystream_a23_source_stride <= 0;
      _mystream_a23_source_sel <= 0;
      _mystream_a23_source_offset_buf <= 0;
      _mystream_a23_source_size_buf <= 0;
      _mystream_a23_source_stride_buf <= 0;
      __variable_wdata_25 <= 0;
      _mystream_a23_source_ram_raddr <= 0;
      _mystream_a23_source_count <= 0;
      _mystream_a24_source_mode <= 5'b0;
      _mystream_a24_source_offset <= 0;
      _mystream_a24_source_size <= 0;
      _mystream_a24_source_stride <= 0;
      _mystream_a24_source_sel <= 0;
      _mystream_a24_source_offset_buf <= 0;
      _mystream_a24_source_size_buf <= 0;
      _mystream_a24_source_stride_buf <= 0;
      __variable_wdata_26 <= 0;
      _mystream_a24_source_ram_raddr <= 0;
      _mystream_a24_source_count <= 0;
      _mystream_a25_source_mode <= 5'b0;
      _mystream_a25_source_offset <= 0;
      _mystream_a25_source_size <= 0;
      _mystream_a25_source_stride <= 0;
      _mystream_a25_source_sel <= 0;
      _mystream_a25_source_offset_buf <= 0;
      _mystream_a25_source_size_buf <= 0;
      _mystream_a25_source_stride_buf <= 0;
      __variable_wdata_27 <= 0;
      _mystream_a25_source_ram_raddr <= 0;
      _mystream_a25_source_count <= 0;
      _mystream_a26_source_mode <= 5'b0;
      _mystream_a26_source_offset <= 0;
      _mystream_a26_source_size <= 0;
      _mystream_a26_source_stride <= 0;
      _mystream_a26_source_sel <= 0;
      _mystream_a26_source_offset_buf <= 0;
      _mystream_a26_source_size_buf <= 0;
      _mystream_a26_source_stride_buf <= 0;
      __variable_wdata_28 <= 0;
      _mystream_a26_source_ram_raddr <= 0;
      _mystream_a26_source_count <= 0;
      _mystream_a27_source_mode <= 5'b0;
      _mystream_a27_source_offset <= 0;
      _mystream_a27_source_size <= 0;
      _mystream_a27_source_stride <= 0;
      _mystream_a27_source_sel <= 0;
      _mystream_a27_source_offset_buf <= 0;
      _mystream_a27_source_size_buf <= 0;
      _mystream_a27_source_stride_buf <= 0;
      __variable_wdata_29 <= 0;
      _mystream_a27_source_ram_raddr <= 0;
      _mystream_a27_source_count <= 0;
      _mystream_a28_source_mode <= 5'b0;
      _mystream_a28_source_offset <= 0;
      _mystream_a28_source_size <= 0;
      _mystream_a28_source_stride <= 0;
      _mystream_a28_source_sel <= 0;
      _mystream_a28_source_offset_buf <= 0;
      _mystream_a28_source_size_buf <= 0;
      _mystream_a28_source_stride_buf <= 0;
      __variable_wdata_30 <= 0;
      _mystream_a28_source_ram_raddr <= 0;
      _mystream_a28_source_count <= 0;
      _mystream_a29_source_mode <= 5'b0;
      _mystream_a29_source_offset <= 0;
      _mystream_a29_source_size <= 0;
      _mystream_a29_source_stride <= 0;
      _mystream_a29_source_sel <= 0;
      _mystream_a29_source_offset_buf <= 0;
      _mystream_a29_source_size_buf <= 0;
      _mystream_a29_source_stride_buf <= 0;
      __variable_wdata_31 <= 0;
      _mystream_a29_source_ram_raddr <= 0;
      _mystream_a29_source_count <= 0;
      _mystream_a30_source_mode <= 5'b0;
      _mystream_a30_source_offset <= 0;
      _mystream_a30_source_size <= 0;
      _mystream_a30_source_stride <= 0;
      _mystream_a30_source_sel <= 0;
      _mystream_a30_source_offset_buf <= 0;
      _mystream_a30_source_size_buf <= 0;
      _mystream_a30_source_stride_buf <= 0;
      __variable_wdata_32 <= 0;
      _mystream_a30_source_ram_raddr <= 0;
      _mystream_a30_source_count <= 0;
      _mystream_a31_source_mode <= 5'b0;
      _mystream_a31_source_offset <= 0;
      _mystream_a31_source_size <= 0;
      _mystream_a31_source_stride <= 0;
      _mystream_a31_source_sel <= 0;
      _mystream_a31_source_offset_buf <= 0;
      _mystream_a31_source_size_buf <= 0;
      _mystream_a31_source_stride_buf <= 0;
      __variable_wdata_33 <= 0;
      _mystream_a31_source_ram_raddr <= 0;
      _mystream_a31_source_count <= 0;
      _mystream_b0_source_mode <= 5'b0;
      _mystream_b0_source_offset <= 0;
      _mystream_b0_source_size <= 0;
      _mystream_b0_source_stride <= 0;
      _mystream_b0_source_sel <= 0;
      _mystream_b0_source_offset_buf <= 0;
      _mystream_b0_source_size_buf <= 0;
      _mystream_b0_source_stride_buf <= 0;
      __variable_wdata_34 <= 0;
      _mystream_b0_source_ram_raddr <= 0;
      _mystream_b0_source_count <= 0;
      _mystream_b1_source_mode <= 5'b0;
      _mystream_b1_source_offset <= 0;
      _mystream_b1_source_size <= 0;
      _mystream_b1_source_stride <= 0;
      _mystream_b1_source_sel <= 0;
      _mystream_b1_source_offset_buf <= 0;
      _mystream_b1_source_size_buf <= 0;
      _mystream_b1_source_stride_buf <= 0;
      __variable_wdata_35 <= 0;
      _mystream_b1_source_ram_raddr <= 0;
      _mystream_b1_source_count <= 0;
      _mystream_b2_source_mode <= 5'b0;
      _mystream_b2_source_offset <= 0;
      _mystream_b2_source_size <= 0;
      _mystream_b2_source_stride <= 0;
      _mystream_b2_source_sel <= 0;
      _mystream_b2_source_offset_buf <= 0;
      _mystream_b2_source_size_buf <= 0;
      _mystream_b2_source_stride_buf <= 0;
      __variable_wdata_36 <= 0;
      _mystream_b2_source_ram_raddr <= 0;
      _mystream_b2_source_count <= 0;
      _mystream_b3_source_mode <= 5'b0;
      _mystream_b3_source_offset <= 0;
      _mystream_b3_source_size <= 0;
      _mystream_b3_source_stride <= 0;
      _mystream_b3_source_sel <= 0;
      _mystream_b3_source_offset_buf <= 0;
      _mystream_b3_source_size_buf <= 0;
      _mystream_b3_source_stride_buf <= 0;
      __variable_wdata_37 <= 0;
      _mystream_b3_source_ram_raddr <= 0;
      _mystream_b3_source_count <= 0;
      _mystream_b4_source_mode <= 5'b0;
      _mystream_b4_source_offset <= 0;
      _mystream_b4_source_size <= 0;
      _mystream_b4_source_stride <= 0;
      _mystream_b4_source_sel <= 0;
      _mystream_b4_source_offset_buf <= 0;
      _mystream_b4_source_size_buf <= 0;
      _mystream_b4_source_stride_buf <= 0;
      __variable_wdata_38 <= 0;
      _mystream_b4_source_ram_raddr <= 0;
      _mystream_b4_source_count <= 0;
      _mystream_b5_source_mode <= 5'b0;
      _mystream_b5_source_offset <= 0;
      _mystream_b5_source_size <= 0;
      _mystream_b5_source_stride <= 0;
      _mystream_b5_source_sel <= 0;
      _mystream_b5_source_offset_buf <= 0;
      _mystream_b5_source_size_buf <= 0;
      _mystream_b5_source_stride_buf <= 0;
      __variable_wdata_39 <= 0;
      _mystream_b5_source_ram_raddr <= 0;
      _mystream_b5_source_count <= 0;
      _mystream_b6_source_mode <= 5'b0;
      _mystream_b6_source_offset <= 0;
      _mystream_b6_source_size <= 0;
      _mystream_b6_source_stride <= 0;
      _mystream_b6_source_sel <= 0;
      _mystream_b6_source_offset_buf <= 0;
      _mystream_b6_source_size_buf <= 0;
      _mystream_b6_source_stride_buf <= 0;
      __variable_wdata_40 <= 0;
      _mystream_b6_source_ram_raddr <= 0;
      _mystream_b6_source_count <= 0;
      _mystream_b7_source_mode <= 5'b0;
      _mystream_b7_source_offset <= 0;
      _mystream_b7_source_size <= 0;
      _mystream_b7_source_stride <= 0;
      _mystream_b7_source_sel <= 0;
      _mystream_b7_source_offset_buf <= 0;
      _mystream_b7_source_size_buf <= 0;
      _mystream_b7_source_stride_buf <= 0;
      __variable_wdata_41 <= 0;
      _mystream_b7_source_ram_raddr <= 0;
      _mystream_b7_source_count <= 0;
      _mystream_b8_source_mode <= 5'b0;
      _mystream_b8_source_offset <= 0;
      _mystream_b8_source_size <= 0;
      _mystream_b8_source_stride <= 0;
      _mystream_b8_source_sel <= 0;
      _mystream_b8_source_offset_buf <= 0;
      _mystream_b8_source_size_buf <= 0;
      _mystream_b8_source_stride_buf <= 0;
      __variable_wdata_42 <= 0;
      _mystream_b8_source_ram_raddr <= 0;
      _mystream_b8_source_count <= 0;
      _mystream_b9_source_mode <= 5'b0;
      _mystream_b9_source_offset <= 0;
      _mystream_b9_source_size <= 0;
      _mystream_b9_source_stride <= 0;
      _mystream_b9_source_sel <= 0;
      _mystream_b9_source_offset_buf <= 0;
      _mystream_b9_source_size_buf <= 0;
      _mystream_b9_source_stride_buf <= 0;
      __variable_wdata_43 <= 0;
      _mystream_b9_source_ram_raddr <= 0;
      _mystream_b9_source_count <= 0;
      _mystream_b10_source_mode <= 5'b0;
      _mystream_b10_source_offset <= 0;
      _mystream_b10_source_size <= 0;
      _mystream_b10_source_stride <= 0;
      _mystream_b10_source_sel <= 0;
      _mystream_b10_source_offset_buf <= 0;
      _mystream_b10_source_size_buf <= 0;
      _mystream_b10_source_stride_buf <= 0;
      __variable_wdata_44 <= 0;
      _mystream_b10_source_ram_raddr <= 0;
      _mystream_b10_source_count <= 0;
      _mystream_b11_source_mode <= 5'b0;
      _mystream_b11_source_offset <= 0;
      _mystream_b11_source_size <= 0;
      _mystream_b11_source_stride <= 0;
      _mystream_b11_source_sel <= 0;
      _mystream_b11_source_offset_buf <= 0;
      _mystream_b11_source_size_buf <= 0;
      _mystream_b11_source_stride_buf <= 0;
      __variable_wdata_45 <= 0;
      _mystream_b11_source_ram_raddr <= 0;
      _mystream_b11_source_count <= 0;
      _mystream_b12_source_mode <= 5'b0;
      _mystream_b12_source_offset <= 0;
      _mystream_b12_source_size <= 0;
      _mystream_b12_source_stride <= 0;
      _mystream_b12_source_sel <= 0;
      _mystream_b12_source_offset_buf <= 0;
      _mystream_b12_source_size_buf <= 0;
      _mystream_b12_source_stride_buf <= 0;
      __variable_wdata_46 <= 0;
      _mystream_b12_source_ram_raddr <= 0;
      _mystream_b12_source_count <= 0;
      _mystream_b13_source_mode <= 5'b0;
      _mystream_b13_source_offset <= 0;
      _mystream_b13_source_size <= 0;
      _mystream_b13_source_stride <= 0;
      _mystream_b13_source_sel <= 0;
      _mystream_b13_source_offset_buf <= 0;
      _mystream_b13_source_size_buf <= 0;
      _mystream_b13_source_stride_buf <= 0;
      __variable_wdata_47 <= 0;
      _mystream_b13_source_ram_raddr <= 0;
      _mystream_b13_source_count <= 0;
      _mystream_b14_source_mode <= 5'b0;
      _mystream_b14_source_offset <= 0;
      _mystream_b14_source_size <= 0;
      _mystream_b14_source_stride <= 0;
      _mystream_b14_source_sel <= 0;
      _mystream_b14_source_offset_buf <= 0;
      _mystream_b14_source_size_buf <= 0;
      _mystream_b14_source_stride_buf <= 0;
      __variable_wdata_48 <= 0;
      _mystream_b14_source_ram_raddr <= 0;
      _mystream_b14_source_count <= 0;
      _mystream_b15_source_mode <= 5'b0;
      _mystream_b15_source_offset <= 0;
      _mystream_b15_source_size <= 0;
      _mystream_b15_source_stride <= 0;
      _mystream_b15_source_sel <= 0;
      _mystream_b15_source_offset_buf <= 0;
      _mystream_b15_source_size_buf <= 0;
      _mystream_b15_source_stride_buf <= 0;
      __variable_wdata_49 <= 0;
      _mystream_b15_source_ram_raddr <= 0;
      _mystream_b15_source_count <= 0;
      _mystream_b16_source_mode <= 5'b0;
      _mystream_b16_source_offset <= 0;
      _mystream_b16_source_size <= 0;
      _mystream_b16_source_stride <= 0;
      _mystream_b16_source_sel <= 0;
      _mystream_b16_source_offset_buf <= 0;
      _mystream_b16_source_size_buf <= 0;
      _mystream_b16_source_stride_buf <= 0;
      __variable_wdata_50 <= 0;
      _mystream_b16_source_ram_raddr <= 0;
      _mystream_b16_source_count <= 0;
      _mystream_b17_source_mode <= 5'b0;
      _mystream_b17_source_offset <= 0;
      _mystream_b17_source_size <= 0;
      _mystream_b17_source_stride <= 0;
      _mystream_b17_source_sel <= 0;
      _mystream_b17_source_offset_buf <= 0;
      _mystream_b17_source_size_buf <= 0;
      _mystream_b17_source_stride_buf <= 0;
      __variable_wdata_51 <= 0;
      _mystream_b17_source_ram_raddr <= 0;
      _mystream_b17_source_count <= 0;
      _mystream_b18_source_mode <= 5'b0;
      _mystream_b18_source_offset <= 0;
      _mystream_b18_source_size <= 0;
      _mystream_b18_source_stride <= 0;
      _mystream_b18_source_sel <= 0;
      _mystream_b18_source_offset_buf <= 0;
      _mystream_b18_source_size_buf <= 0;
      _mystream_b18_source_stride_buf <= 0;
      __variable_wdata_52 <= 0;
      _mystream_b18_source_ram_raddr <= 0;
      _mystream_b18_source_count <= 0;
      _mystream_b19_source_mode <= 5'b0;
      _mystream_b19_source_offset <= 0;
      _mystream_b19_source_size <= 0;
      _mystream_b19_source_stride <= 0;
      _mystream_b19_source_sel <= 0;
      _mystream_b19_source_offset_buf <= 0;
      _mystream_b19_source_size_buf <= 0;
      _mystream_b19_source_stride_buf <= 0;
      __variable_wdata_53 <= 0;
      _mystream_b19_source_ram_raddr <= 0;
      _mystream_b19_source_count <= 0;
      _mystream_b20_source_mode <= 5'b0;
      _mystream_b20_source_offset <= 0;
      _mystream_b20_source_size <= 0;
      _mystream_b20_source_stride <= 0;
      _mystream_b20_source_sel <= 0;
      _mystream_b20_source_offset_buf <= 0;
      _mystream_b20_source_size_buf <= 0;
      _mystream_b20_source_stride_buf <= 0;
      __variable_wdata_54 <= 0;
      _mystream_b20_source_ram_raddr <= 0;
      _mystream_b20_source_count <= 0;
      _mystream_b21_source_mode <= 5'b0;
      _mystream_b21_source_offset <= 0;
      _mystream_b21_source_size <= 0;
      _mystream_b21_source_stride <= 0;
      _mystream_b21_source_sel <= 0;
      _mystream_b21_source_offset_buf <= 0;
      _mystream_b21_source_size_buf <= 0;
      _mystream_b21_source_stride_buf <= 0;
      __variable_wdata_55 <= 0;
      _mystream_b21_source_ram_raddr <= 0;
      _mystream_b21_source_count <= 0;
      _mystream_b22_source_mode <= 5'b0;
      _mystream_b22_source_offset <= 0;
      _mystream_b22_source_size <= 0;
      _mystream_b22_source_stride <= 0;
      _mystream_b22_source_sel <= 0;
      _mystream_b22_source_offset_buf <= 0;
      _mystream_b22_source_size_buf <= 0;
      _mystream_b22_source_stride_buf <= 0;
      __variable_wdata_56 <= 0;
      _mystream_b22_source_ram_raddr <= 0;
      _mystream_b22_source_count <= 0;
      _mystream_b23_source_mode <= 5'b0;
      _mystream_b23_source_offset <= 0;
      _mystream_b23_source_size <= 0;
      _mystream_b23_source_stride <= 0;
      _mystream_b23_source_sel <= 0;
      _mystream_b23_source_offset_buf <= 0;
      _mystream_b23_source_size_buf <= 0;
      _mystream_b23_source_stride_buf <= 0;
      __variable_wdata_57 <= 0;
      _mystream_b23_source_ram_raddr <= 0;
      _mystream_b23_source_count <= 0;
      _mystream_b24_source_mode <= 5'b0;
      _mystream_b24_source_offset <= 0;
      _mystream_b24_source_size <= 0;
      _mystream_b24_source_stride <= 0;
      _mystream_b24_source_sel <= 0;
      _mystream_b24_source_offset_buf <= 0;
      _mystream_b24_source_size_buf <= 0;
      _mystream_b24_source_stride_buf <= 0;
      __variable_wdata_58 <= 0;
      _mystream_b24_source_ram_raddr <= 0;
      _mystream_b24_source_count <= 0;
      _mystream_b25_source_mode <= 5'b0;
      _mystream_b25_source_offset <= 0;
      _mystream_b25_source_size <= 0;
      _mystream_b25_source_stride <= 0;
      _mystream_b25_source_sel <= 0;
      _mystream_b25_source_offset_buf <= 0;
      _mystream_b25_source_size_buf <= 0;
      _mystream_b25_source_stride_buf <= 0;
      __variable_wdata_59 <= 0;
      _mystream_b25_source_ram_raddr <= 0;
      _mystream_b25_source_count <= 0;
      _mystream_b26_source_mode <= 5'b0;
      _mystream_b26_source_offset <= 0;
      _mystream_b26_source_size <= 0;
      _mystream_b26_source_stride <= 0;
      _mystream_b26_source_sel <= 0;
      _mystream_b26_source_offset_buf <= 0;
      _mystream_b26_source_size_buf <= 0;
      _mystream_b26_source_stride_buf <= 0;
      __variable_wdata_60 <= 0;
      _mystream_b26_source_ram_raddr <= 0;
      _mystream_b26_source_count <= 0;
      _mystream_b27_source_mode <= 5'b0;
      _mystream_b27_source_offset <= 0;
      _mystream_b27_source_size <= 0;
      _mystream_b27_source_stride <= 0;
      _mystream_b27_source_sel <= 0;
      _mystream_b27_source_offset_buf <= 0;
      _mystream_b27_source_size_buf <= 0;
      _mystream_b27_source_stride_buf <= 0;
      __variable_wdata_61 <= 0;
      _mystream_b27_source_ram_raddr <= 0;
      _mystream_b27_source_count <= 0;
      _mystream_b28_source_mode <= 5'b0;
      _mystream_b28_source_offset <= 0;
      _mystream_b28_source_size <= 0;
      _mystream_b28_source_stride <= 0;
      _mystream_b28_source_sel <= 0;
      _mystream_b28_source_offset_buf <= 0;
      _mystream_b28_source_size_buf <= 0;
      _mystream_b28_source_stride_buf <= 0;
      __variable_wdata_62 <= 0;
      _mystream_b28_source_ram_raddr <= 0;
      _mystream_b28_source_count <= 0;
      _mystream_b29_source_mode <= 5'b0;
      _mystream_b29_source_offset <= 0;
      _mystream_b29_source_size <= 0;
      _mystream_b29_source_stride <= 0;
      _mystream_b29_source_sel <= 0;
      _mystream_b29_source_offset_buf <= 0;
      _mystream_b29_source_size_buf <= 0;
      _mystream_b29_source_stride_buf <= 0;
      __variable_wdata_63 <= 0;
      _mystream_b29_source_ram_raddr <= 0;
      _mystream_b29_source_count <= 0;
      _mystream_b30_source_mode <= 5'b0;
      _mystream_b30_source_offset <= 0;
      _mystream_b30_source_size <= 0;
      _mystream_b30_source_stride <= 0;
      _mystream_b30_source_sel <= 0;
      _mystream_b30_source_offset_buf <= 0;
      _mystream_b30_source_size_buf <= 0;
      _mystream_b30_source_stride_buf <= 0;
      __variable_wdata_64 <= 0;
      _mystream_b30_source_ram_raddr <= 0;
      _mystream_b30_source_count <= 0;
      _mystream_b31_source_mode <= 5'b0;
      _mystream_b31_source_offset <= 0;
      _mystream_b31_source_size <= 0;
      _mystream_b31_source_stride <= 0;
      _mystream_b31_source_sel <= 0;
      _mystream_b31_source_offset_buf <= 0;
      _mystream_b31_source_size_buf <= 0;
      _mystream_b31_source_stride_buf <= 0;
      __variable_wdata_65 <= 0;
      _mystream_b31_source_ram_raddr <= 0;
      _mystream_b31_source_count <= 0;
      _tmp_378 <= 0;
      _tmp_379 <= 0;
      _tmp_380 <= 0;
      _tmp_381 <= 0;
      _tmp_382 <= 0;
      _tmp_383 <= 0;
      _tmp_384 <= 0;
      _tmp_385 <= 0;
      _tmp_386 <= 0;
      _tmp_387 <= 0;
      _tmp_388 <= 0;
      _tmp_389 <= 0;
      _tmp_392 <= 0;
      _tmp_393 <= 0;
      _tmp_394 <= 0;
      _tmp_395 <= 0;
      _tmp_396 <= 0;
      _tmp_397 <= 0;
      _mystream_sum_vec0_sink_mode <= 5'b0;
      _mystream_sum_vec0_sink_offset <= 0;
      _mystream_sum_vec0_sink_size <= 0;
      _mystream_sum_vec0_sink_stride <= 0;
      _mystream_sum_vec0_sink_sel <= 0;
      _mystream_sum_vec0_sink_offset_buf <= 0;
      _mystream_sum_vec0_sink_size_buf <= 0;
      _mystream_sum_vec0_sink_stride_buf <= 0;
      _mystream_sum_vec0_sink_waddr <= 0;
      _mystream_sum_vec0_sink_count <= 0;
      _mystream_sum_vec0_sink_wdata <= 0;
      _tmp_399 <= 0;
      _tmp_400 <= 0;
      _tmp_401 <= 0;
      _tmp_402 <= 0;
      _tmp_403 <= 0;
      _tmp_404 <= 0;
      _tmp_405 <= 0;
      _tmp_406 <= 0;
      _tmp_407 <= 0;
      _tmp_408 <= 0;
      _tmp_409 <= 0;
      _tmp_410 <= 0;
      _tmp_413 <= 0;
      _tmp_414 <= 0;
      _tmp_415 <= 0;
      _tmp_416 <= 0;
      _tmp_417 <= 0;
      _tmp_418 <= 0;
      _mystream_sum_vec1_sink_mode <= 5'b0;
      _mystream_sum_vec1_sink_offset <= 0;
      _mystream_sum_vec1_sink_size <= 0;
      _mystream_sum_vec1_sink_stride <= 0;
      _mystream_sum_vec1_sink_sel <= 0;
      _mystream_sum_vec1_sink_offset_buf <= 0;
      _mystream_sum_vec1_sink_size_buf <= 0;
      _mystream_sum_vec1_sink_stride_buf <= 0;
      _mystream_sum_vec1_sink_waddr <= 0;
      _mystream_sum_vec1_sink_count <= 0;
      _mystream_sum_vec1_sink_wdata <= 0;
      _tmp_420 <= 0;
      _tmp_421 <= 0;
      _tmp_422 <= 0;
      _tmp_423 <= 0;
      _tmp_424 <= 0;
      _tmp_425 <= 0;
      _tmp_426 <= 0;
      _tmp_427 <= 0;
      _tmp_428 <= 0;
      _tmp_429 <= 0;
      _tmp_430 <= 0;
      _tmp_431 <= 0;
      _tmp_434 <= 0;
      _tmp_435 <= 0;
      _tmp_436 <= 0;
      _tmp_437 <= 0;
      _tmp_438 <= 0;
      _tmp_439 <= 0;
      _mystream_sum_vec2_sink_mode <= 5'b0;
      _mystream_sum_vec2_sink_offset <= 0;
      _mystream_sum_vec2_sink_size <= 0;
      _mystream_sum_vec2_sink_stride <= 0;
      _mystream_sum_vec2_sink_sel <= 0;
      _mystream_sum_vec2_sink_offset_buf <= 0;
      _mystream_sum_vec2_sink_size_buf <= 0;
      _mystream_sum_vec2_sink_stride_buf <= 0;
      _mystream_sum_vec2_sink_waddr <= 0;
      _mystream_sum_vec2_sink_count <= 0;
      _mystream_sum_vec2_sink_wdata <= 0;
      _tmp_441 <= 0;
      _tmp_442 <= 0;
      _tmp_443 <= 0;
      _tmp_444 <= 0;
      _tmp_445 <= 0;
      _tmp_446 <= 0;
      _tmp_447 <= 0;
      _tmp_448 <= 0;
      _tmp_449 <= 0;
      _tmp_450 <= 0;
      _tmp_451 <= 0;
      _tmp_452 <= 0;
      _tmp_455 <= 0;
      _tmp_456 <= 0;
      _tmp_457 <= 0;
      _tmp_458 <= 0;
      _tmp_459 <= 0;
      _tmp_460 <= 0;
      _mystream_sum_vec3_sink_mode <= 5'b0;
      _mystream_sum_vec3_sink_offset <= 0;
      _mystream_sum_vec3_sink_size <= 0;
      _mystream_sum_vec3_sink_stride <= 0;
      _mystream_sum_vec3_sink_sel <= 0;
      _mystream_sum_vec3_sink_offset_buf <= 0;
      _mystream_sum_vec3_sink_size_buf <= 0;
      _mystream_sum_vec3_sink_stride_buf <= 0;
      _mystream_sum_vec3_sink_waddr <= 0;
      _mystream_sum_vec3_sink_count <= 0;
      _mystream_sum_vec3_sink_wdata <= 0;
      _tmp_462 <= 0;
      _tmp_463 <= 0;
      _tmp_464 <= 0;
      _tmp_465 <= 0;
      _tmp_466 <= 0;
      _tmp_467 <= 0;
      _tmp_468 <= 0;
      _tmp_469 <= 0;
      _tmp_470 <= 0;
      _tmp_471 <= 0;
      _tmp_472 <= 0;
      _tmp_473 <= 0;
      _tmp_476 <= 0;
      _tmp_477 <= 0;
      _tmp_478 <= 0;
      _tmp_479 <= 0;
      _tmp_480 <= 0;
      _tmp_481 <= 0;
      _mystream_sum_vec4_sink_mode <= 5'b0;
      _mystream_sum_vec4_sink_offset <= 0;
      _mystream_sum_vec4_sink_size <= 0;
      _mystream_sum_vec4_sink_stride <= 0;
      _mystream_sum_vec4_sink_sel <= 0;
      _mystream_sum_vec4_sink_offset_buf <= 0;
      _mystream_sum_vec4_sink_size_buf <= 0;
      _mystream_sum_vec4_sink_stride_buf <= 0;
      _mystream_sum_vec4_sink_waddr <= 0;
      _mystream_sum_vec4_sink_count <= 0;
      _mystream_sum_vec4_sink_wdata <= 0;
      _tmp_483 <= 0;
      _tmp_484 <= 0;
      _tmp_485 <= 0;
      _tmp_486 <= 0;
      _tmp_487 <= 0;
      _tmp_488 <= 0;
      _tmp_489 <= 0;
      _tmp_490 <= 0;
      _tmp_491 <= 0;
      _tmp_492 <= 0;
      _tmp_493 <= 0;
      _tmp_494 <= 0;
      _tmp_497 <= 0;
      _tmp_498 <= 0;
      _tmp_499 <= 0;
      _tmp_500 <= 0;
      _tmp_501 <= 0;
      _tmp_502 <= 0;
      _mystream_sum_vec5_sink_mode <= 5'b0;
      _mystream_sum_vec5_sink_offset <= 0;
      _mystream_sum_vec5_sink_size <= 0;
      _mystream_sum_vec5_sink_stride <= 0;
      _mystream_sum_vec5_sink_sel <= 0;
      _mystream_sum_vec5_sink_offset_buf <= 0;
      _mystream_sum_vec5_sink_size_buf <= 0;
      _mystream_sum_vec5_sink_stride_buf <= 0;
      _mystream_sum_vec5_sink_waddr <= 0;
      _mystream_sum_vec5_sink_count <= 0;
      _mystream_sum_vec5_sink_wdata <= 0;
      _tmp_504 <= 0;
      _tmp_505 <= 0;
      _tmp_506 <= 0;
      _tmp_507 <= 0;
      _tmp_508 <= 0;
      _tmp_509 <= 0;
      _tmp_510 <= 0;
      _tmp_511 <= 0;
      _tmp_512 <= 0;
      _tmp_513 <= 0;
      _tmp_514 <= 0;
      _tmp_515 <= 0;
      _tmp_518 <= 0;
      _tmp_519 <= 0;
      _tmp_520 <= 0;
      _tmp_521 <= 0;
      _tmp_522 <= 0;
      _tmp_523 <= 0;
      _mystream_sum_vec6_sink_mode <= 5'b0;
      _mystream_sum_vec6_sink_offset <= 0;
      _mystream_sum_vec6_sink_size <= 0;
      _mystream_sum_vec6_sink_stride <= 0;
      _mystream_sum_vec6_sink_sel <= 0;
      _mystream_sum_vec6_sink_offset_buf <= 0;
      _mystream_sum_vec6_sink_size_buf <= 0;
      _mystream_sum_vec6_sink_stride_buf <= 0;
      _mystream_sum_vec6_sink_waddr <= 0;
      _mystream_sum_vec6_sink_count <= 0;
      _mystream_sum_vec6_sink_wdata <= 0;
      _tmp_525 <= 0;
      _tmp_526 <= 0;
      _tmp_527 <= 0;
      _tmp_528 <= 0;
      _tmp_529 <= 0;
      _tmp_530 <= 0;
      _tmp_531 <= 0;
      _tmp_532 <= 0;
      _tmp_533 <= 0;
      _tmp_534 <= 0;
      _tmp_535 <= 0;
      _tmp_536 <= 0;
      _tmp_539 <= 0;
      _tmp_540 <= 0;
      _tmp_541 <= 0;
      _tmp_542 <= 0;
      _tmp_543 <= 0;
      _tmp_544 <= 0;
      _mystream_sum_vec7_sink_mode <= 5'b0;
      _mystream_sum_vec7_sink_offset <= 0;
      _mystream_sum_vec7_sink_size <= 0;
      _mystream_sum_vec7_sink_stride <= 0;
      _mystream_sum_vec7_sink_sel <= 0;
      _mystream_sum_vec7_sink_offset_buf <= 0;
      _mystream_sum_vec7_sink_size_buf <= 0;
      _mystream_sum_vec7_sink_stride_buf <= 0;
      _mystream_sum_vec7_sink_waddr <= 0;
      _mystream_sum_vec7_sink_count <= 0;
      _mystream_sum_vec7_sink_wdata <= 0;
      _tmp_546 <= 0;
      _tmp_547 <= 0;
      _tmp_548 <= 0;
      _tmp_549 <= 0;
      _tmp_550 <= 0;
      _tmp_551 <= 0;
      _tmp_552 <= 0;
      _tmp_553 <= 0;
      _tmp_554 <= 0;
      _tmp_555 <= 0;
      _tmp_556 <= 0;
      _tmp_557 <= 0;
      _tmp_560 <= 0;
      _tmp_561 <= 0;
      _tmp_562 <= 0;
      _tmp_563 <= 0;
      _tmp_564 <= 0;
      _tmp_565 <= 0;
      _mystream_sum_vec8_sink_mode <= 5'b0;
      _mystream_sum_vec8_sink_offset <= 0;
      _mystream_sum_vec8_sink_size <= 0;
      _mystream_sum_vec8_sink_stride <= 0;
      _mystream_sum_vec8_sink_sel <= 0;
      _mystream_sum_vec8_sink_offset_buf <= 0;
      _mystream_sum_vec8_sink_size_buf <= 0;
      _mystream_sum_vec8_sink_stride_buf <= 0;
      _mystream_sum_vec8_sink_waddr <= 0;
      _mystream_sum_vec8_sink_count <= 0;
      _mystream_sum_vec8_sink_wdata <= 0;
      _tmp_567 <= 0;
      _tmp_568 <= 0;
      _tmp_569 <= 0;
      _tmp_570 <= 0;
      _tmp_571 <= 0;
      _tmp_572 <= 0;
      _tmp_573 <= 0;
      _tmp_574 <= 0;
      _tmp_575 <= 0;
      _tmp_576 <= 0;
      _tmp_577 <= 0;
      _tmp_578 <= 0;
      _tmp_581 <= 0;
      _tmp_582 <= 0;
      _tmp_583 <= 0;
      _tmp_584 <= 0;
      _tmp_585 <= 0;
      _tmp_586 <= 0;
      _mystream_sum_vec9_sink_mode <= 5'b0;
      _mystream_sum_vec9_sink_offset <= 0;
      _mystream_sum_vec9_sink_size <= 0;
      _mystream_sum_vec9_sink_stride <= 0;
      _mystream_sum_vec9_sink_sel <= 0;
      _mystream_sum_vec9_sink_offset_buf <= 0;
      _mystream_sum_vec9_sink_size_buf <= 0;
      _mystream_sum_vec9_sink_stride_buf <= 0;
      _mystream_sum_vec9_sink_waddr <= 0;
      _mystream_sum_vec9_sink_count <= 0;
      _mystream_sum_vec9_sink_wdata <= 0;
      _tmp_588 <= 0;
      _tmp_589 <= 0;
      _tmp_590 <= 0;
      _tmp_591 <= 0;
      _tmp_592 <= 0;
      _tmp_593 <= 0;
      _tmp_594 <= 0;
      _tmp_595 <= 0;
      _tmp_596 <= 0;
      _tmp_597 <= 0;
      _tmp_598 <= 0;
      _tmp_599 <= 0;
      _tmp_602 <= 0;
      _tmp_603 <= 0;
      _tmp_604 <= 0;
      _tmp_605 <= 0;
      _tmp_606 <= 0;
      _tmp_607 <= 0;
      _mystream_sum_vec10_sink_mode <= 5'b0;
      _mystream_sum_vec10_sink_offset <= 0;
      _mystream_sum_vec10_sink_size <= 0;
      _mystream_sum_vec10_sink_stride <= 0;
      _mystream_sum_vec10_sink_sel <= 0;
      _mystream_sum_vec10_sink_offset_buf <= 0;
      _mystream_sum_vec10_sink_size_buf <= 0;
      _mystream_sum_vec10_sink_stride_buf <= 0;
      _mystream_sum_vec10_sink_waddr <= 0;
      _mystream_sum_vec10_sink_count <= 0;
      _mystream_sum_vec10_sink_wdata <= 0;
      _tmp_609 <= 0;
      _tmp_610 <= 0;
      _tmp_611 <= 0;
      _tmp_612 <= 0;
      _tmp_613 <= 0;
      _tmp_614 <= 0;
      _tmp_615 <= 0;
      _tmp_616 <= 0;
      _tmp_617 <= 0;
      _tmp_618 <= 0;
      _tmp_619 <= 0;
      _tmp_620 <= 0;
      _tmp_623 <= 0;
      _tmp_624 <= 0;
      _tmp_625 <= 0;
      _tmp_626 <= 0;
      _tmp_627 <= 0;
      _tmp_628 <= 0;
      _mystream_sum_vec11_sink_mode <= 5'b0;
      _mystream_sum_vec11_sink_offset <= 0;
      _mystream_sum_vec11_sink_size <= 0;
      _mystream_sum_vec11_sink_stride <= 0;
      _mystream_sum_vec11_sink_sel <= 0;
      _mystream_sum_vec11_sink_offset_buf <= 0;
      _mystream_sum_vec11_sink_size_buf <= 0;
      _mystream_sum_vec11_sink_stride_buf <= 0;
      _mystream_sum_vec11_sink_waddr <= 0;
      _mystream_sum_vec11_sink_count <= 0;
      _mystream_sum_vec11_sink_wdata <= 0;
      _tmp_630 <= 0;
      _tmp_631 <= 0;
      _tmp_632 <= 0;
      _tmp_633 <= 0;
      _tmp_634 <= 0;
      _tmp_635 <= 0;
      _tmp_636 <= 0;
      _tmp_637 <= 0;
      _tmp_638 <= 0;
      _tmp_639 <= 0;
      _tmp_640 <= 0;
      _tmp_641 <= 0;
      _tmp_644 <= 0;
      _tmp_645 <= 0;
      _tmp_646 <= 0;
      _tmp_647 <= 0;
      _tmp_648 <= 0;
      _tmp_649 <= 0;
      _mystream_sum_vec12_sink_mode <= 5'b0;
      _mystream_sum_vec12_sink_offset <= 0;
      _mystream_sum_vec12_sink_size <= 0;
      _mystream_sum_vec12_sink_stride <= 0;
      _mystream_sum_vec12_sink_sel <= 0;
      _mystream_sum_vec12_sink_offset_buf <= 0;
      _mystream_sum_vec12_sink_size_buf <= 0;
      _mystream_sum_vec12_sink_stride_buf <= 0;
      _mystream_sum_vec12_sink_waddr <= 0;
      _mystream_sum_vec12_sink_count <= 0;
      _mystream_sum_vec12_sink_wdata <= 0;
      _tmp_651 <= 0;
      _tmp_652 <= 0;
      _tmp_653 <= 0;
      _tmp_654 <= 0;
      _tmp_655 <= 0;
      _tmp_656 <= 0;
      _tmp_657 <= 0;
      _tmp_658 <= 0;
      _tmp_659 <= 0;
      _tmp_660 <= 0;
      _tmp_661 <= 0;
      _tmp_662 <= 0;
      _tmp_665 <= 0;
      _tmp_666 <= 0;
      _tmp_667 <= 0;
      _tmp_668 <= 0;
      _tmp_669 <= 0;
      _tmp_670 <= 0;
      _mystream_sum_vec13_sink_mode <= 5'b0;
      _mystream_sum_vec13_sink_offset <= 0;
      _mystream_sum_vec13_sink_size <= 0;
      _mystream_sum_vec13_sink_stride <= 0;
      _mystream_sum_vec13_sink_sel <= 0;
      _mystream_sum_vec13_sink_offset_buf <= 0;
      _mystream_sum_vec13_sink_size_buf <= 0;
      _mystream_sum_vec13_sink_stride_buf <= 0;
      _mystream_sum_vec13_sink_waddr <= 0;
      _mystream_sum_vec13_sink_count <= 0;
      _mystream_sum_vec13_sink_wdata <= 0;
      _tmp_672 <= 0;
      _tmp_673 <= 0;
      _tmp_674 <= 0;
      _tmp_675 <= 0;
      _tmp_676 <= 0;
      _tmp_677 <= 0;
      _tmp_678 <= 0;
      _tmp_679 <= 0;
      _tmp_680 <= 0;
      _tmp_681 <= 0;
      _tmp_682 <= 0;
      _tmp_683 <= 0;
      _tmp_686 <= 0;
      _tmp_687 <= 0;
      _tmp_688 <= 0;
      _tmp_689 <= 0;
      _tmp_690 <= 0;
      _tmp_691 <= 0;
      _mystream_sum_vec14_sink_mode <= 5'b0;
      _mystream_sum_vec14_sink_offset <= 0;
      _mystream_sum_vec14_sink_size <= 0;
      _mystream_sum_vec14_sink_stride <= 0;
      _mystream_sum_vec14_sink_sel <= 0;
      _mystream_sum_vec14_sink_offset_buf <= 0;
      _mystream_sum_vec14_sink_size_buf <= 0;
      _mystream_sum_vec14_sink_stride_buf <= 0;
      _mystream_sum_vec14_sink_waddr <= 0;
      _mystream_sum_vec14_sink_count <= 0;
      _mystream_sum_vec14_sink_wdata <= 0;
      _tmp_693 <= 0;
      _tmp_694 <= 0;
      _tmp_695 <= 0;
      _tmp_696 <= 0;
      _tmp_697 <= 0;
      _tmp_698 <= 0;
      _tmp_699 <= 0;
      _tmp_700 <= 0;
      _tmp_701 <= 0;
      _tmp_702 <= 0;
      _tmp_703 <= 0;
      _tmp_704 <= 0;
      _tmp_707 <= 0;
      _tmp_708 <= 0;
      _tmp_709 <= 0;
      _tmp_710 <= 0;
      _tmp_711 <= 0;
      _tmp_712 <= 0;
      _mystream_sum_vec15_sink_mode <= 5'b0;
      _mystream_sum_vec15_sink_offset <= 0;
      _mystream_sum_vec15_sink_size <= 0;
      _mystream_sum_vec15_sink_stride <= 0;
      _mystream_sum_vec15_sink_sel <= 0;
      _mystream_sum_vec15_sink_offset_buf <= 0;
      _mystream_sum_vec15_sink_size_buf <= 0;
      _mystream_sum_vec15_sink_stride_buf <= 0;
      _mystream_sum_vec15_sink_waddr <= 0;
      _mystream_sum_vec15_sink_count <= 0;
      _mystream_sum_vec15_sink_wdata <= 0;
      _tmp_714 <= 0;
      _tmp_715 <= 0;
      _tmp_716 <= 0;
      _tmp_717 <= 0;
      _tmp_718 <= 0;
      _tmp_719 <= 0;
      _tmp_720 <= 0;
      _tmp_721 <= 0;
      _tmp_722 <= 0;
      _tmp_723 <= 0;
      _tmp_724 <= 0;
      _tmp_725 <= 0;
      _tmp_728 <= 0;
      _tmp_729 <= 0;
      _tmp_730 <= 0;
      _tmp_731 <= 0;
      _tmp_732 <= 0;
      _tmp_733 <= 0;
      _mystream_sum_vec16_sink_mode <= 5'b0;
      _mystream_sum_vec16_sink_offset <= 0;
      _mystream_sum_vec16_sink_size <= 0;
      _mystream_sum_vec16_sink_stride <= 0;
      _mystream_sum_vec16_sink_sel <= 0;
      _mystream_sum_vec16_sink_offset_buf <= 0;
      _mystream_sum_vec16_sink_size_buf <= 0;
      _mystream_sum_vec16_sink_stride_buf <= 0;
      _mystream_sum_vec16_sink_waddr <= 0;
      _mystream_sum_vec16_sink_count <= 0;
      _mystream_sum_vec16_sink_wdata <= 0;
      _tmp_735 <= 0;
      _tmp_736 <= 0;
      _tmp_737 <= 0;
      _tmp_738 <= 0;
      _tmp_739 <= 0;
      _tmp_740 <= 0;
      _tmp_741 <= 0;
      _tmp_742 <= 0;
      _tmp_743 <= 0;
      _tmp_744 <= 0;
      _tmp_745 <= 0;
      _tmp_746 <= 0;
      _tmp_749 <= 0;
      _tmp_750 <= 0;
      _tmp_751 <= 0;
      _tmp_752 <= 0;
      _tmp_753 <= 0;
      _tmp_754 <= 0;
      _mystream_sum_vec17_sink_mode <= 5'b0;
      _mystream_sum_vec17_sink_offset <= 0;
      _mystream_sum_vec17_sink_size <= 0;
      _mystream_sum_vec17_sink_stride <= 0;
      _mystream_sum_vec17_sink_sel <= 0;
      _mystream_sum_vec17_sink_offset_buf <= 0;
      _mystream_sum_vec17_sink_size_buf <= 0;
      _mystream_sum_vec17_sink_stride_buf <= 0;
      _mystream_sum_vec17_sink_waddr <= 0;
      _mystream_sum_vec17_sink_count <= 0;
      _mystream_sum_vec17_sink_wdata <= 0;
      _tmp_756 <= 0;
      _tmp_757 <= 0;
      _tmp_758 <= 0;
      _tmp_759 <= 0;
      _tmp_760 <= 0;
      _tmp_761 <= 0;
      _tmp_762 <= 0;
      _tmp_763 <= 0;
      _tmp_764 <= 0;
      _tmp_765 <= 0;
      _tmp_766 <= 0;
      _tmp_767 <= 0;
      _tmp_770 <= 0;
      _tmp_771 <= 0;
      _tmp_772 <= 0;
      _tmp_773 <= 0;
      _tmp_774 <= 0;
      _tmp_775 <= 0;
      _mystream_sum_vec18_sink_mode <= 5'b0;
      _mystream_sum_vec18_sink_offset <= 0;
      _mystream_sum_vec18_sink_size <= 0;
      _mystream_sum_vec18_sink_stride <= 0;
      _mystream_sum_vec18_sink_sel <= 0;
      _mystream_sum_vec18_sink_offset_buf <= 0;
      _mystream_sum_vec18_sink_size_buf <= 0;
      _mystream_sum_vec18_sink_stride_buf <= 0;
      _mystream_sum_vec18_sink_waddr <= 0;
      _mystream_sum_vec18_sink_count <= 0;
      _mystream_sum_vec18_sink_wdata <= 0;
      _tmp_777 <= 0;
      _tmp_778 <= 0;
      _tmp_779 <= 0;
      _tmp_780 <= 0;
      _tmp_781 <= 0;
      _tmp_782 <= 0;
      _tmp_783 <= 0;
      _tmp_784 <= 0;
      _tmp_785 <= 0;
      _tmp_786 <= 0;
      _tmp_787 <= 0;
      _tmp_788 <= 0;
      _tmp_791 <= 0;
      _tmp_792 <= 0;
      _tmp_793 <= 0;
      _tmp_794 <= 0;
      _tmp_795 <= 0;
      _tmp_796 <= 0;
      _mystream_sum_vec19_sink_mode <= 5'b0;
      _mystream_sum_vec19_sink_offset <= 0;
      _mystream_sum_vec19_sink_size <= 0;
      _mystream_sum_vec19_sink_stride <= 0;
      _mystream_sum_vec19_sink_sel <= 0;
      _mystream_sum_vec19_sink_offset_buf <= 0;
      _mystream_sum_vec19_sink_size_buf <= 0;
      _mystream_sum_vec19_sink_stride_buf <= 0;
      _mystream_sum_vec19_sink_waddr <= 0;
      _mystream_sum_vec19_sink_count <= 0;
      _mystream_sum_vec19_sink_wdata <= 0;
      _tmp_798 <= 0;
      _tmp_799 <= 0;
      _tmp_800 <= 0;
      _tmp_801 <= 0;
      _tmp_802 <= 0;
      _tmp_803 <= 0;
      _tmp_804 <= 0;
      _tmp_805 <= 0;
      _tmp_806 <= 0;
      _tmp_807 <= 0;
      _tmp_808 <= 0;
      _tmp_809 <= 0;
      _tmp_812 <= 0;
      _tmp_813 <= 0;
      _tmp_814 <= 0;
      _tmp_815 <= 0;
      _tmp_816 <= 0;
      _tmp_817 <= 0;
      _mystream_sum_vec20_sink_mode <= 5'b0;
      _mystream_sum_vec20_sink_offset <= 0;
      _mystream_sum_vec20_sink_size <= 0;
      _mystream_sum_vec20_sink_stride <= 0;
      _mystream_sum_vec20_sink_sel <= 0;
      _mystream_sum_vec20_sink_offset_buf <= 0;
      _mystream_sum_vec20_sink_size_buf <= 0;
      _mystream_sum_vec20_sink_stride_buf <= 0;
      _mystream_sum_vec20_sink_waddr <= 0;
      _mystream_sum_vec20_sink_count <= 0;
      _mystream_sum_vec20_sink_wdata <= 0;
      _tmp_819 <= 0;
      _tmp_820 <= 0;
      _tmp_821 <= 0;
      _tmp_822 <= 0;
      _tmp_823 <= 0;
      _tmp_824 <= 0;
      _tmp_825 <= 0;
      _tmp_826 <= 0;
      _tmp_827 <= 0;
      _tmp_828 <= 0;
      _tmp_829 <= 0;
      _tmp_830 <= 0;
      _tmp_833 <= 0;
      _tmp_834 <= 0;
      _tmp_835 <= 0;
      _tmp_836 <= 0;
      _tmp_837 <= 0;
      _tmp_838 <= 0;
      _mystream_sum_vec21_sink_mode <= 5'b0;
      _mystream_sum_vec21_sink_offset <= 0;
      _mystream_sum_vec21_sink_size <= 0;
      _mystream_sum_vec21_sink_stride <= 0;
      _mystream_sum_vec21_sink_sel <= 0;
      _mystream_sum_vec21_sink_offset_buf <= 0;
      _mystream_sum_vec21_sink_size_buf <= 0;
      _mystream_sum_vec21_sink_stride_buf <= 0;
      _mystream_sum_vec21_sink_waddr <= 0;
      _mystream_sum_vec21_sink_count <= 0;
      _mystream_sum_vec21_sink_wdata <= 0;
      _tmp_840 <= 0;
      _tmp_841 <= 0;
      _tmp_842 <= 0;
      _tmp_843 <= 0;
      _tmp_844 <= 0;
      _tmp_845 <= 0;
      _tmp_846 <= 0;
      _tmp_847 <= 0;
      _tmp_848 <= 0;
      _tmp_849 <= 0;
      _tmp_850 <= 0;
      _tmp_851 <= 0;
      _tmp_854 <= 0;
      _tmp_855 <= 0;
      _tmp_856 <= 0;
      _tmp_857 <= 0;
      _tmp_858 <= 0;
      _tmp_859 <= 0;
      _mystream_sum_vec22_sink_mode <= 5'b0;
      _mystream_sum_vec22_sink_offset <= 0;
      _mystream_sum_vec22_sink_size <= 0;
      _mystream_sum_vec22_sink_stride <= 0;
      _mystream_sum_vec22_sink_sel <= 0;
      _mystream_sum_vec22_sink_offset_buf <= 0;
      _mystream_sum_vec22_sink_size_buf <= 0;
      _mystream_sum_vec22_sink_stride_buf <= 0;
      _mystream_sum_vec22_sink_waddr <= 0;
      _mystream_sum_vec22_sink_count <= 0;
      _mystream_sum_vec22_sink_wdata <= 0;
      _tmp_861 <= 0;
      _tmp_862 <= 0;
      _tmp_863 <= 0;
      _tmp_864 <= 0;
      _tmp_865 <= 0;
      _tmp_866 <= 0;
      _tmp_867 <= 0;
      _tmp_868 <= 0;
      _tmp_869 <= 0;
      _tmp_870 <= 0;
      _tmp_871 <= 0;
      _tmp_872 <= 0;
      _tmp_875 <= 0;
      _tmp_876 <= 0;
      _tmp_877 <= 0;
      _tmp_878 <= 0;
      _tmp_879 <= 0;
      _tmp_880 <= 0;
      _mystream_sum_vec23_sink_mode <= 5'b0;
      _mystream_sum_vec23_sink_offset <= 0;
      _mystream_sum_vec23_sink_size <= 0;
      _mystream_sum_vec23_sink_stride <= 0;
      _mystream_sum_vec23_sink_sel <= 0;
      _mystream_sum_vec23_sink_offset_buf <= 0;
      _mystream_sum_vec23_sink_size_buf <= 0;
      _mystream_sum_vec23_sink_stride_buf <= 0;
      _mystream_sum_vec23_sink_waddr <= 0;
      _mystream_sum_vec23_sink_count <= 0;
      _mystream_sum_vec23_sink_wdata <= 0;
      _tmp_882 <= 0;
      _tmp_883 <= 0;
      _tmp_884 <= 0;
      _tmp_885 <= 0;
      _tmp_886 <= 0;
      _tmp_887 <= 0;
      _tmp_888 <= 0;
      _tmp_889 <= 0;
      _tmp_890 <= 0;
      _tmp_891 <= 0;
      _tmp_892 <= 0;
      _tmp_893 <= 0;
      _tmp_896 <= 0;
      _tmp_897 <= 0;
      _tmp_898 <= 0;
      _tmp_899 <= 0;
      _tmp_900 <= 0;
      _tmp_901 <= 0;
      _mystream_sum_vec24_sink_mode <= 5'b0;
      _mystream_sum_vec24_sink_offset <= 0;
      _mystream_sum_vec24_sink_size <= 0;
      _mystream_sum_vec24_sink_stride <= 0;
      _mystream_sum_vec24_sink_sel <= 0;
      _mystream_sum_vec24_sink_offset_buf <= 0;
      _mystream_sum_vec24_sink_size_buf <= 0;
      _mystream_sum_vec24_sink_stride_buf <= 0;
      _mystream_sum_vec24_sink_waddr <= 0;
      _mystream_sum_vec24_sink_count <= 0;
      _mystream_sum_vec24_sink_wdata <= 0;
      _tmp_903 <= 0;
      _tmp_904 <= 0;
      _tmp_905 <= 0;
      _tmp_906 <= 0;
      _tmp_907 <= 0;
      _tmp_908 <= 0;
      _tmp_909 <= 0;
      _tmp_910 <= 0;
      _tmp_911 <= 0;
      _tmp_912 <= 0;
      _tmp_913 <= 0;
      _tmp_914 <= 0;
      _tmp_917 <= 0;
      _tmp_918 <= 0;
      _tmp_919 <= 0;
      _tmp_920 <= 0;
      _tmp_921 <= 0;
      _tmp_922 <= 0;
      _mystream_sum_vec25_sink_mode <= 5'b0;
      _mystream_sum_vec25_sink_offset <= 0;
      _mystream_sum_vec25_sink_size <= 0;
      _mystream_sum_vec25_sink_stride <= 0;
      _mystream_sum_vec25_sink_sel <= 0;
      _mystream_sum_vec25_sink_offset_buf <= 0;
      _mystream_sum_vec25_sink_size_buf <= 0;
      _mystream_sum_vec25_sink_stride_buf <= 0;
      _mystream_sum_vec25_sink_waddr <= 0;
      _mystream_sum_vec25_sink_count <= 0;
      _mystream_sum_vec25_sink_wdata <= 0;
      _tmp_924 <= 0;
      _tmp_925 <= 0;
      _tmp_926 <= 0;
      _tmp_927 <= 0;
      _tmp_928 <= 0;
      _tmp_929 <= 0;
      _tmp_930 <= 0;
      _tmp_931 <= 0;
      _tmp_932 <= 0;
      _tmp_933 <= 0;
      _tmp_934 <= 0;
      _tmp_935 <= 0;
      _tmp_938 <= 0;
      _tmp_939 <= 0;
      _tmp_940 <= 0;
      _tmp_941 <= 0;
      _tmp_942 <= 0;
      _tmp_943 <= 0;
      _mystream_sum_vec26_sink_mode <= 5'b0;
      _mystream_sum_vec26_sink_offset <= 0;
      _mystream_sum_vec26_sink_size <= 0;
      _mystream_sum_vec26_sink_stride <= 0;
      _mystream_sum_vec26_sink_sel <= 0;
      _mystream_sum_vec26_sink_offset_buf <= 0;
      _mystream_sum_vec26_sink_size_buf <= 0;
      _mystream_sum_vec26_sink_stride_buf <= 0;
      _mystream_sum_vec26_sink_waddr <= 0;
      _mystream_sum_vec26_sink_count <= 0;
      _mystream_sum_vec26_sink_wdata <= 0;
      _tmp_945 <= 0;
      _tmp_946 <= 0;
      _tmp_947 <= 0;
      _tmp_948 <= 0;
      _tmp_949 <= 0;
      _tmp_950 <= 0;
      _tmp_951 <= 0;
      _tmp_952 <= 0;
      _tmp_953 <= 0;
      _tmp_954 <= 0;
      _tmp_955 <= 0;
      _tmp_956 <= 0;
      _tmp_959 <= 0;
      _tmp_960 <= 0;
      _tmp_961 <= 0;
      _tmp_962 <= 0;
      _tmp_963 <= 0;
      _tmp_964 <= 0;
      _mystream_sum_vec27_sink_mode <= 5'b0;
      _mystream_sum_vec27_sink_offset <= 0;
      _mystream_sum_vec27_sink_size <= 0;
      _mystream_sum_vec27_sink_stride <= 0;
      _mystream_sum_vec27_sink_sel <= 0;
      _mystream_sum_vec27_sink_offset_buf <= 0;
      _mystream_sum_vec27_sink_size_buf <= 0;
      _mystream_sum_vec27_sink_stride_buf <= 0;
      _mystream_sum_vec27_sink_waddr <= 0;
      _mystream_sum_vec27_sink_count <= 0;
      _mystream_sum_vec27_sink_wdata <= 0;
      _tmp_966 <= 0;
      _tmp_967 <= 0;
      _tmp_968 <= 0;
      _tmp_969 <= 0;
      _tmp_970 <= 0;
      _tmp_971 <= 0;
      _tmp_972 <= 0;
      _tmp_973 <= 0;
      _tmp_974 <= 0;
      _tmp_975 <= 0;
      _tmp_976 <= 0;
      _tmp_977 <= 0;
      _tmp_980 <= 0;
      _tmp_981 <= 0;
      _tmp_982 <= 0;
      _tmp_983 <= 0;
      _tmp_984 <= 0;
      _tmp_985 <= 0;
      _mystream_sum_vec28_sink_mode <= 5'b0;
      _mystream_sum_vec28_sink_offset <= 0;
      _mystream_sum_vec28_sink_size <= 0;
      _mystream_sum_vec28_sink_stride <= 0;
      _mystream_sum_vec28_sink_sel <= 0;
      _mystream_sum_vec28_sink_offset_buf <= 0;
      _mystream_sum_vec28_sink_size_buf <= 0;
      _mystream_sum_vec28_sink_stride_buf <= 0;
      _mystream_sum_vec28_sink_waddr <= 0;
      _mystream_sum_vec28_sink_count <= 0;
      _mystream_sum_vec28_sink_wdata <= 0;
      _tmp_987 <= 0;
      _tmp_988 <= 0;
      _tmp_989 <= 0;
      _tmp_990 <= 0;
      _tmp_991 <= 0;
      _tmp_992 <= 0;
      _tmp_993 <= 0;
      _tmp_994 <= 0;
      _tmp_995 <= 0;
      _tmp_996 <= 0;
      _tmp_997 <= 0;
      _tmp_998 <= 0;
      _tmp_1001 <= 0;
      _tmp_1002 <= 0;
      _tmp_1003 <= 0;
      _tmp_1004 <= 0;
      _tmp_1005 <= 0;
      _tmp_1006 <= 0;
      _mystream_sum_vec29_sink_mode <= 5'b0;
      _mystream_sum_vec29_sink_offset <= 0;
      _mystream_sum_vec29_sink_size <= 0;
      _mystream_sum_vec29_sink_stride <= 0;
      _mystream_sum_vec29_sink_sel <= 0;
      _mystream_sum_vec29_sink_offset_buf <= 0;
      _mystream_sum_vec29_sink_size_buf <= 0;
      _mystream_sum_vec29_sink_stride_buf <= 0;
      _mystream_sum_vec29_sink_waddr <= 0;
      _mystream_sum_vec29_sink_count <= 0;
      _mystream_sum_vec29_sink_wdata <= 0;
      _tmp_1008 <= 0;
      _tmp_1009 <= 0;
      _tmp_1010 <= 0;
      _tmp_1011 <= 0;
      _tmp_1012 <= 0;
      _tmp_1013 <= 0;
      _tmp_1014 <= 0;
      _tmp_1015 <= 0;
      _tmp_1016 <= 0;
      _tmp_1017 <= 0;
      _tmp_1018 <= 0;
      _tmp_1019 <= 0;
      _tmp_1022 <= 0;
      _tmp_1023 <= 0;
      _tmp_1024 <= 0;
      _tmp_1025 <= 0;
      _tmp_1026 <= 0;
      _tmp_1027 <= 0;
      _mystream_sum_vec30_sink_mode <= 5'b0;
      _mystream_sum_vec30_sink_offset <= 0;
      _mystream_sum_vec30_sink_size <= 0;
      _mystream_sum_vec30_sink_stride <= 0;
      _mystream_sum_vec30_sink_sel <= 0;
      _mystream_sum_vec30_sink_offset_buf <= 0;
      _mystream_sum_vec30_sink_size_buf <= 0;
      _mystream_sum_vec30_sink_stride_buf <= 0;
      _mystream_sum_vec30_sink_waddr <= 0;
      _mystream_sum_vec30_sink_count <= 0;
      _mystream_sum_vec30_sink_wdata <= 0;
      _tmp_1029 <= 0;
      _tmp_1030 <= 0;
      _tmp_1031 <= 0;
      _tmp_1032 <= 0;
      _tmp_1033 <= 0;
      _tmp_1034 <= 0;
      _tmp_1035 <= 0;
      _tmp_1036 <= 0;
      _tmp_1037 <= 0;
      _tmp_1038 <= 0;
      _tmp_1039 <= 0;
      _tmp_1040 <= 0;
      _tmp_1043 <= 0;
      _tmp_1044 <= 0;
      _tmp_1045 <= 0;
      _tmp_1046 <= 0;
      _tmp_1047 <= 0;
      _tmp_1048 <= 0;
      _mystream_sum_vec31_sink_mode <= 5'b0;
      _mystream_sum_vec31_sink_offset <= 0;
      _mystream_sum_vec31_sink_size <= 0;
      _mystream_sum_vec31_sink_stride <= 0;
      _mystream_sum_vec31_sink_sel <= 0;
      _mystream_sum_vec31_sink_offset_buf <= 0;
      _mystream_sum_vec31_sink_size_buf <= 0;
      _mystream_sum_vec31_sink_stride_buf <= 0;
      _mystream_sum_vec31_sink_waddr <= 0;
      _mystream_sum_vec31_sink_count <= 0;
      _mystream_sum_vec31_sink_wdata <= 0;
      _tmp_1050 <= 0;
      _tmp_1051 <= 0;
      _tmp_1052 <= 0;
      _tmp_1053 <= 0;
      _tmp_1054 <= 0;
      _tmp_1055 <= 0;
      __variable_wdata_130 <= 0;
      _tmp_1056 <= 0;
      _tmp_1057 <= 0;
      _tmp_1058 <= 0;
      _tmp_1059 <= 0;
      _tmp_1062 <= 0;
      _tmp_1065 <= 0;
      _tmp_1066 <= 0;
      _tmp_1067 <= 0;
      _tmp_1068 <= 0;
      _tmp_1069 <= 0;
      _tmp_1070 <= 0;
      _tmp_1071 <= 0;
      _tmp_1072 <= 0;
      _tmp_1073 <= 0;
      _tmp_1074 <= 0;
      _tmp_1075 <= 0;
      _tmp_1076 <= 0;
      _tmp_1077 <= 0;
      _tmp_1078 <= 0;
      _tmp_1079 <= 0;
      _tmp_1080 <= 0;
      _tmp_1081 <= 0;
      _tmp_1082 <= 0;
      _tmp_1083 <= 0;
      _tmp_1084 <= 0;
      _mystream_busy_reg <= 0;
    end else begin
      if(_mystream_stream_oready) begin
        _mystream_a0_source_ram_renable <= 0;
        _mystream_a0_source_fifo_deq <= 0;
      end 
      _mystream_a0_idle <= _mystream_a0_idle;
      if(_mystream_stream_oready) begin
        _mystream_a1_source_ram_renable <= 0;
        _mystream_a1_source_fifo_deq <= 0;
      end 
      _mystream_a1_idle <= _mystream_a1_idle;
      if(_mystream_stream_oready) begin
        _mystream_a2_source_ram_renable <= 0;
        _mystream_a2_source_fifo_deq <= 0;
      end 
      _mystream_a2_idle <= _mystream_a2_idle;
      if(_mystream_stream_oready) begin
        _mystream_a3_source_ram_renable <= 0;
        _mystream_a3_source_fifo_deq <= 0;
      end 
      _mystream_a3_idle <= _mystream_a3_idle;
      if(_mystream_stream_oready) begin
        _mystream_a4_source_ram_renable <= 0;
        _mystream_a4_source_fifo_deq <= 0;
      end 
      _mystream_a4_idle <= _mystream_a4_idle;
      if(_mystream_stream_oready) begin
        _mystream_a5_source_ram_renable <= 0;
        _mystream_a5_source_fifo_deq <= 0;
      end 
      _mystream_a5_idle <= _mystream_a5_idle;
      if(_mystream_stream_oready) begin
        _mystream_a6_source_ram_renable <= 0;
        _mystream_a6_source_fifo_deq <= 0;
      end 
      _mystream_a6_idle <= _mystream_a6_idle;
      if(_mystream_stream_oready) begin
        _mystream_a7_source_ram_renable <= 0;
        _mystream_a7_source_fifo_deq <= 0;
      end 
      _mystream_a7_idle <= _mystream_a7_idle;
      if(_mystream_stream_oready) begin
        _mystream_a8_source_ram_renable <= 0;
        _mystream_a8_source_fifo_deq <= 0;
      end 
      _mystream_a8_idle <= _mystream_a8_idle;
      if(_mystream_stream_oready) begin
        _mystream_a9_source_ram_renable <= 0;
        _mystream_a9_source_fifo_deq <= 0;
      end 
      _mystream_a9_idle <= _mystream_a9_idle;
      if(_mystream_stream_oready) begin
        _mystream_a10_source_ram_renable <= 0;
        _mystream_a10_source_fifo_deq <= 0;
      end 
      _mystream_a10_idle <= _mystream_a10_idle;
      if(_mystream_stream_oready) begin
        _mystream_a11_source_ram_renable <= 0;
        _mystream_a11_source_fifo_deq <= 0;
      end 
      _mystream_a11_idle <= _mystream_a11_idle;
      if(_mystream_stream_oready) begin
        _mystream_a12_source_ram_renable <= 0;
        _mystream_a12_source_fifo_deq <= 0;
      end 
      _mystream_a12_idle <= _mystream_a12_idle;
      if(_mystream_stream_oready) begin
        _mystream_a13_source_ram_renable <= 0;
        _mystream_a13_source_fifo_deq <= 0;
      end 
      _mystream_a13_idle <= _mystream_a13_idle;
      if(_mystream_stream_oready) begin
        _mystream_a14_source_ram_renable <= 0;
        _mystream_a14_source_fifo_deq <= 0;
      end 
      _mystream_a14_idle <= _mystream_a14_idle;
      if(_mystream_stream_oready) begin
        _mystream_a15_source_ram_renable <= 0;
        _mystream_a15_source_fifo_deq <= 0;
      end 
      _mystream_a15_idle <= _mystream_a15_idle;
      if(_mystream_stream_oready) begin
        _mystream_a16_source_ram_renable <= 0;
        _mystream_a16_source_fifo_deq <= 0;
      end 
      _mystream_a16_idle <= _mystream_a16_idle;
      if(_mystream_stream_oready) begin
        _mystream_a17_source_ram_renable <= 0;
        _mystream_a17_source_fifo_deq <= 0;
      end 
      _mystream_a17_idle <= _mystream_a17_idle;
      if(_mystream_stream_oready) begin
        _mystream_a18_source_ram_renable <= 0;
        _mystream_a18_source_fifo_deq <= 0;
      end 
      _mystream_a18_idle <= _mystream_a18_idle;
      if(_mystream_stream_oready) begin
        _mystream_a19_source_ram_renable <= 0;
        _mystream_a19_source_fifo_deq <= 0;
      end 
      _mystream_a19_idle <= _mystream_a19_idle;
      if(_mystream_stream_oready) begin
        _mystream_a20_source_ram_renable <= 0;
        _mystream_a20_source_fifo_deq <= 0;
      end 
      _mystream_a20_idle <= _mystream_a20_idle;
      if(_mystream_stream_oready) begin
        _mystream_a21_source_ram_renable <= 0;
        _mystream_a21_source_fifo_deq <= 0;
      end 
      _mystream_a21_idle <= _mystream_a21_idle;
      if(_mystream_stream_oready) begin
        _mystream_a22_source_ram_renable <= 0;
        _mystream_a22_source_fifo_deq <= 0;
      end 
      _mystream_a22_idle <= _mystream_a22_idle;
      if(_mystream_stream_oready) begin
        _mystream_a23_source_ram_renable <= 0;
        _mystream_a23_source_fifo_deq <= 0;
      end 
      _mystream_a23_idle <= _mystream_a23_idle;
      if(_mystream_stream_oready) begin
        _mystream_a24_source_ram_renable <= 0;
        _mystream_a24_source_fifo_deq <= 0;
      end 
      _mystream_a24_idle <= _mystream_a24_idle;
      if(_mystream_stream_oready) begin
        _mystream_a25_source_ram_renable <= 0;
        _mystream_a25_source_fifo_deq <= 0;
      end 
      _mystream_a25_idle <= _mystream_a25_idle;
      if(_mystream_stream_oready) begin
        _mystream_a26_source_ram_renable <= 0;
        _mystream_a26_source_fifo_deq <= 0;
      end 
      _mystream_a26_idle <= _mystream_a26_idle;
      if(_mystream_stream_oready) begin
        _mystream_a27_source_ram_renable <= 0;
        _mystream_a27_source_fifo_deq <= 0;
      end 
      _mystream_a27_idle <= _mystream_a27_idle;
      if(_mystream_stream_oready) begin
        _mystream_a28_source_ram_renable <= 0;
        _mystream_a28_source_fifo_deq <= 0;
      end 
      _mystream_a28_idle <= _mystream_a28_idle;
      if(_mystream_stream_oready) begin
        _mystream_a29_source_ram_renable <= 0;
        _mystream_a29_source_fifo_deq <= 0;
      end 
      _mystream_a29_idle <= _mystream_a29_idle;
      if(_mystream_stream_oready) begin
        _mystream_a30_source_ram_renable <= 0;
        _mystream_a30_source_fifo_deq <= 0;
      end 
      _mystream_a30_idle <= _mystream_a30_idle;
      if(_mystream_stream_oready) begin
        _mystream_a31_source_ram_renable <= 0;
        _mystream_a31_source_fifo_deq <= 0;
      end 
      _mystream_a31_idle <= _mystream_a31_idle;
      if(_mystream_stream_oready) begin
        _mystream_b0_source_ram_renable <= 0;
        _mystream_b0_source_fifo_deq <= 0;
      end 
      _mystream_b0_idle <= _mystream_b0_idle;
      if(_mystream_stream_oready) begin
        _mystream_b1_source_ram_renable <= 0;
        _mystream_b1_source_fifo_deq <= 0;
      end 
      _mystream_b1_idle <= _mystream_b1_idle;
      if(_mystream_stream_oready) begin
        _mystream_b2_source_ram_renable <= 0;
        _mystream_b2_source_fifo_deq <= 0;
      end 
      _mystream_b2_idle <= _mystream_b2_idle;
      if(_mystream_stream_oready) begin
        _mystream_b3_source_ram_renable <= 0;
        _mystream_b3_source_fifo_deq <= 0;
      end 
      _mystream_b3_idle <= _mystream_b3_idle;
      if(_mystream_stream_oready) begin
        _mystream_b4_source_ram_renable <= 0;
        _mystream_b4_source_fifo_deq <= 0;
      end 
      _mystream_b4_idle <= _mystream_b4_idle;
      if(_mystream_stream_oready) begin
        _mystream_b5_source_ram_renable <= 0;
        _mystream_b5_source_fifo_deq <= 0;
      end 
      _mystream_b5_idle <= _mystream_b5_idle;
      if(_mystream_stream_oready) begin
        _mystream_b6_source_ram_renable <= 0;
        _mystream_b6_source_fifo_deq <= 0;
      end 
      _mystream_b6_idle <= _mystream_b6_idle;
      if(_mystream_stream_oready) begin
        _mystream_b7_source_ram_renable <= 0;
        _mystream_b7_source_fifo_deq <= 0;
      end 
      _mystream_b7_idle <= _mystream_b7_idle;
      if(_mystream_stream_oready) begin
        _mystream_b8_source_ram_renable <= 0;
        _mystream_b8_source_fifo_deq <= 0;
      end 
      _mystream_b8_idle <= _mystream_b8_idle;
      if(_mystream_stream_oready) begin
        _mystream_b9_source_ram_renable <= 0;
        _mystream_b9_source_fifo_deq <= 0;
      end 
      _mystream_b9_idle <= _mystream_b9_idle;
      if(_mystream_stream_oready) begin
        _mystream_b10_source_ram_renable <= 0;
        _mystream_b10_source_fifo_deq <= 0;
      end 
      _mystream_b10_idle <= _mystream_b10_idle;
      if(_mystream_stream_oready) begin
        _mystream_b11_source_ram_renable <= 0;
        _mystream_b11_source_fifo_deq <= 0;
      end 
      _mystream_b11_idle <= _mystream_b11_idle;
      if(_mystream_stream_oready) begin
        _mystream_b12_source_ram_renable <= 0;
        _mystream_b12_source_fifo_deq <= 0;
      end 
      _mystream_b12_idle <= _mystream_b12_idle;
      if(_mystream_stream_oready) begin
        _mystream_b13_source_ram_renable <= 0;
        _mystream_b13_source_fifo_deq <= 0;
      end 
      _mystream_b13_idle <= _mystream_b13_idle;
      if(_mystream_stream_oready) begin
        _mystream_b14_source_ram_renable <= 0;
        _mystream_b14_source_fifo_deq <= 0;
      end 
      _mystream_b14_idle <= _mystream_b14_idle;
      if(_mystream_stream_oready) begin
        _mystream_b15_source_ram_renable <= 0;
        _mystream_b15_source_fifo_deq <= 0;
      end 
      _mystream_b15_idle <= _mystream_b15_idle;
      if(_mystream_stream_oready) begin
        _mystream_b16_source_ram_renable <= 0;
        _mystream_b16_source_fifo_deq <= 0;
      end 
      _mystream_b16_idle <= _mystream_b16_idle;
      if(_mystream_stream_oready) begin
        _mystream_b17_source_ram_renable <= 0;
        _mystream_b17_source_fifo_deq <= 0;
      end 
      _mystream_b17_idle <= _mystream_b17_idle;
      if(_mystream_stream_oready) begin
        _mystream_b18_source_ram_renable <= 0;
        _mystream_b18_source_fifo_deq <= 0;
      end 
      _mystream_b18_idle <= _mystream_b18_idle;
      if(_mystream_stream_oready) begin
        _mystream_b19_source_ram_renable <= 0;
        _mystream_b19_source_fifo_deq <= 0;
      end 
      _mystream_b19_idle <= _mystream_b19_idle;
      if(_mystream_stream_oready) begin
        _mystream_b20_source_ram_renable <= 0;
        _mystream_b20_source_fifo_deq <= 0;
      end 
      _mystream_b20_idle <= _mystream_b20_idle;
      if(_mystream_stream_oready) begin
        _mystream_b21_source_ram_renable <= 0;
        _mystream_b21_source_fifo_deq <= 0;
      end 
      _mystream_b21_idle <= _mystream_b21_idle;
      if(_mystream_stream_oready) begin
        _mystream_b22_source_ram_renable <= 0;
        _mystream_b22_source_fifo_deq <= 0;
      end 
      _mystream_b22_idle <= _mystream_b22_idle;
      if(_mystream_stream_oready) begin
        _mystream_b23_source_ram_renable <= 0;
        _mystream_b23_source_fifo_deq <= 0;
      end 
      _mystream_b23_idle <= _mystream_b23_idle;
      if(_mystream_stream_oready) begin
        _mystream_b24_source_ram_renable <= 0;
        _mystream_b24_source_fifo_deq <= 0;
      end 
      _mystream_b24_idle <= _mystream_b24_idle;
      if(_mystream_stream_oready) begin
        _mystream_b25_source_ram_renable <= 0;
        _mystream_b25_source_fifo_deq <= 0;
      end 
      _mystream_b25_idle <= _mystream_b25_idle;
      if(_mystream_stream_oready) begin
        _mystream_b26_source_ram_renable <= 0;
        _mystream_b26_source_fifo_deq <= 0;
      end 
      _mystream_b26_idle <= _mystream_b26_idle;
      if(_mystream_stream_oready) begin
        _mystream_b27_source_ram_renable <= 0;
        _mystream_b27_source_fifo_deq <= 0;
      end 
      _mystream_b27_idle <= _mystream_b27_idle;
      if(_mystream_stream_oready) begin
        _mystream_b28_source_ram_renable <= 0;
        _mystream_b28_source_fifo_deq <= 0;
      end 
      _mystream_b28_idle <= _mystream_b28_idle;
      if(_mystream_stream_oready) begin
        _mystream_b29_source_ram_renable <= 0;
        _mystream_b29_source_fifo_deq <= 0;
      end 
      _mystream_b29_idle <= _mystream_b29_idle;
      if(_mystream_stream_oready) begin
        _mystream_b30_source_ram_renable <= 0;
        _mystream_b30_source_fifo_deq <= 0;
      end 
      _mystream_b30_idle <= _mystream_b30_idle;
      if(_mystream_stream_oready) begin
        _mystream_b31_source_ram_renable <= 0;
        _mystream_b31_source_fifo_deq <= 0;
      end 
      _mystream_b31_idle <= _mystream_b31_idle;
      if(_mystream_stream_oready) begin
        _mystream_bias0_source_ram_renable <= 0;
        _mystream_bias0_source_fifo_deq <= 0;
      end 
      _mystream_bias0_idle <= _mystream_bias0_idle;
      if(_mystream_stream_oready) begin
        _mystream_bias1_source_ram_renable <= 0;
        _mystream_bias1_source_fifo_deq <= 0;
      end 
      _mystream_bias1_idle <= _mystream_bias1_idle;
      if(_mystream_stream_oready) begin
        _mystream_bias2_source_ram_renable <= 0;
        _mystream_bias2_source_fifo_deq <= 0;
      end 
      _mystream_bias2_idle <= _mystream_bias2_idle;
      if(_mystream_stream_oready) begin
        _mystream_bias3_source_ram_renable <= 0;
        _mystream_bias3_source_fifo_deq <= 0;
      end 
      _mystream_bias3_idle <= _mystream_bias3_idle;
      if(_mystream_stream_oready) begin
        _mystream_bias4_source_ram_renable <= 0;
        _mystream_bias4_source_fifo_deq <= 0;
      end 
      _mystream_bias4_idle <= _mystream_bias4_idle;
      if(_mystream_stream_oready) begin
        _mystream_bias5_source_ram_renable <= 0;
        _mystream_bias5_source_fifo_deq <= 0;
      end 
      _mystream_bias5_idle <= _mystream_bias5_idle;
      if(_mystream_stream_oready) begin
        _mystream_bias6_source_ram_renable <= 0;
        _mystream_bias6_source_fifo_deq <= 0;
      end 
      _mystream_bias6_idle <= _mystream_bias6_idle;
      if(_mystream_stream_oready) begin
        _mystream_bias7_source_ram_renable <= 0;
        _mystream_bias7_source_fifo_deq <= 0;
      end 
      _mystream_bias7_idle <= _mystream_bias7_idle;
      if(_mystream_stream_oready) begin
        _mystream_bias8_source_ram_renable <= 0;
        _mystream_bias8_source_fifo_deq <= 0;
      end 
      _mystream_bias8_idle <= _mystream_bias8_idle;
      if(_mystream_stream_oready) begin
        _mystream_bias9_source_ram_renable <= 0;
        _mystream_bias9_source_fifo_deq <= 0;
      end 
      _mystream_bias9_idle <= _mystream_bias9_idle;
      if(_mystream_stream_oready) begin
        _mystream_bias10_source_ram_renable <= 0;
        _mystream_bias10_source_fifo_deq <= 0;
      end 
      _mystream_bias10_idle <= _mystream_bias10_idle;
      if(_mystream_stream_oready) begin
        _mystream_bias11_source_ram_renable <= 0;
        _mystream_bias11_source_fifo_deq <= 0;
      end 
      _mystream_bias11_idle <= _mystream_bias11_idle;
      if(_mystream_stream_oready) begin
        _mystream_bias12_source_ram_renable <= 0;
        _mystream_bias12_source_fifo_deq <= 0;
      end 
      _mystream_bias12_idle <= _mystream_bias12_idle;
      if(_mystream_stream_oready) begin
        _mystream_bias13_source_ram_renable <= 0;
        _mystream_bias13_source_fifo_deq <= 0;
      end 
      _mystream_bias13_idle <= _mystream_bias13_idle;
      if(_mystream_stream_oready) begin
        _mystream_bias14_source_ram_renable <= 0;
        _mystream_bias14_source_fifo_deq <= 0;
      end 
      _mystream_bias14_idle <= _mystream_bias14_idle;
      if(_mystream_stream_oready) begin
        _mystream_bias15_source_ram_renable <= 0;
        _mystream_bias15_source_fifo_deq <= 0;
      end 
      _mystream_bias15_idle <= _mystream_bias15_idle;
      if(_mystream_stream_oready) begin
        _mystream_bias16_source_ram_renable <= 0;
        _mystream_bias16_source_fifo_deq <= 0;
      end 
      _mystream_bias16_idle <= _mystream_bias16_idle;
      if(_mystream_stream_oready) begin
        _mystream_bias17_source_ram_renable <= 0;
        _mystream_bias17_source_fifo_deq <= 0;
      end 
      _mystream_bias17_idle <= _mystream_bias17_idle;
      if(_mystream_stream_oready) begin
        _mystream_bias18_source_ram_renable <= 0;
        _mystream_bias18_source_fifo_deq <= 0;
      end 
      _mystream_bias18_idle <= _mystream_bias18_idle;
      if(_mystream_stream_oready) begin
        _mystream_bias19_source_ram_renable <= 0;
        _mystream_bias19_source_fifo_deq <= 0;
      end 
      _mystream_bias19_idle <= _mystream_bias19_idle;
      if(_mystream_stream_oready) begin
        _mystream_bias20_source_ram_renable <= 0;
        _mystream_bias20_source_fifo_deq <= 0;
      end 
      _mystream_bias20_idle <= _mystream_bias20_idle;
      if(_mystream_stream_oready) begin
        _mystream_bias21_source_ram_renable <= 0;
        _mystream_bias21_source_fifo_deq <= 0;
      end 
      _mystream_bias21_idle <= _mystream_bias21_idle;
      if(_mystream_stream_oready) begin
        _mystream_bias22_source_ram_renable <= 0;
        _mystream_bias22_source_fifo_deq <= 0;
      end 
      _mystream_bias22_idle <= _mystream_bias22_idle;
      if(_mystream_stream_oready) begin
        _mystream_bias23_source_ram_renable <= 0;
        _mystream_bias23_source_fifo_deq <= 0;
      end 
      _mystream_bias23_idle <= _mystream_bias23_idle;
      if(_mystream_stream_oready) begin
        _mystream_bias24_source_ram_renable <= 0;
        _mystream_bias24_source_fifo_deq <= 0;
      end 
      _mystream_bias24_idle <= _mystream_bias24_idle;
      if(_mystream_stream_oready) begin
        _mystream_bias25_source_ram_renable <= 0;
        _mystream_bias25_source_fifo_deq <= 0;
      end 
      _mystream_bias25_idle <= _mystream_bias25_idle;
      if(_mystream_stream_oready) begin
        _mystream_bias26_source_ram_renable <= 0;
        _mystream_bias26_source_fifo_deq <= 0;
      end 
      _mystream_bias26_idle <= _mystream_bias26_idle;
      if(_mystream_stream_oready) begin
        _mystream_bias27_source_ram_renable <= 0;
        _mystream_bias27_source_fifo_deq <= 0;
      end 
      _mystream_bias27_idle <= _mystream_bias27_idle;
      if(_mystream_stream_oready) begin
        _mystream_bias28_source_ram_renable <= 0;
        _mystream_bias28_source_fifo_deq <= 0;
      end 
      _mystream_bias28_idle <= _mystream_bias28_idle;
      if(_mystream_stream_oready) begin
        _mystream_bias29_source_ram_renable <= 0;
        _mystream_bias29_source_fifo_deq <= 0;
      end 
      _mystream_bias29_idle <= _mystream_bias29_idle;
      if(_mystream_stream_oready) begin
        _mystream_bias30_source_ram_renable <= 0;
        _mystream_bias30_source_fifo_deq <= 0;
      end 
      _mystream_bias30_idle <= _mystream_bias30_idle;
      if(_mystream_stream_oready) begin
        _mystream_bias31_source_ram_renable <= 0;
        _mystream_bias31_source_fifo_deq <= 0;
      end 
      _mystream_bias31_idle <= _mystream_bias31_idle;
      if(_mystream_stream_oready) begin
        _mystream_sum_vec0_sink_wenable <= 0;
        _mystream_sum_vec0_sink_fifo_enq <= 0;
      end 
      if(_mystream_stream_oready) begin
        _mystream_sum_vec1_sink_wenable <= 0;
        _mystream_sum_vec1_sink_fifo_enq <= 0;
      end 
      if(_mystream_stream_oready) begin
        _mystream_sum_vec2_sink_wenable <= 0;
        _mystream_sum_vec2_sink_fifo_enq <= 0;
      end 
      if(_mystream_stream_oready) begin
        _mystream_sum_vec3_sink_wenable <= 0;
        _mystream_sum_vec3_sink_fifo_enq <= 0;
      end 
      if(_mystream_stream_oready) begin
        _mystream_sum_vec4_sink_wenable <= 0;
        _mystream_sum_vec4_sink_fifo_enq <= 0;
      end 
      if(_mystream_stream_oready) begin
        _mystream_sum_vec5_sink_wenable <= 0;
        _mystream_sum_vec5_sink_fifo_enq <= 0;
      end 
      if(_mystream_stream_oready) begin
        _mystream_sum_vec6_sink_wenable <= 0;
        _mystream_sum_vec6_sink_fifo_enq <= 0;
      end 
      if(_mystream_stream_oready) begin
        _mystream_sum_vec7_sink_wenable <= 0;
        _mystream_sum_vec7_sink_fifo_enq <= 0;
      end 
      if(_mystream_stream_oready) begin
        _mystream_sum_vec8_sink_wenable <= 0;
        _mystream_sum_vec8_sink_fifo_enq <= 0;
      end 
      if(_mystream_stream_oready) begin
        _mystream_sum_vec9_sink_wenable <= 0;
        _mystream_sum_vec9_sink_fifo_enq <= 0;
      end 
      if(_mystream_stream_oready) begin
        _mystream_sum_vec10_sink_wenable <= 0;
        _mystream_sum_vec10_sink_fifo_enq <= 0;
      end 
      if(_mystream_stream_oready) begin
        _mystream_sum_vec11_sink_wenable <= 0;
        _mystream_sum_vec11_sink_fifo_enq <= 0;
      end 
      if(_mystream_stream_oready) begin
        _mystream_sum_vec12_sink_wenable <= 0;
        _mystream_sum_vec12_sink_fifo_enq <= 0;
      end 
      if(_mystream_stream_oready) begin
        _mystream_sum_vec13_sink_wenable <= 0;
        _mystream_sum_vec13_sink_fifo_enq <= 0;
      end 
      if(_mystream_stream_oready) begin
        _mystream_sum_vec14_sink_wenable <= 0;
        _mystream_sum_vec14_sink_fifo_enq <= 0;
      end 
      if(_mystream_stream_oready) begin
        _mystream_sum_vec15_sink_wenable <= 0;
        _mystream_sum_vec15_sink_fifo_enq <= 0;
      end 
      if(_mystream_stream_oready) begin
        _mystream_sum_vec16_sink_wenable <= 0;
        _mystream_sum_vec16_sink_fifo_enq <= 0;
      end 
      if(_mystream_stream_oready) begin
        _mystream_sum_vec17_sink_wenable <= 0;
        _mystream_sum_vec17_sink_fifo_enq <= 0;
      end 
      if(_mystream_stream_oready) begin
        _mystream_sum_vec18_sink_wenable <= 0;
        _mystream_sum_vec18_sink_fifo_enq <= 0;
      end 
      if(_mystream_stream_oready) begin
        _mystream_sum_vec19_sink_wenable <= 0;
        _mystream_sum_vec19_sink_fifo_enq <= 0;
      end 
      if(_mystream_stream_oready) begin
        _mystream_sum_vec20_sink_wenable <= 0;
        _mystream_sum_vec20_sink_fifo_enq <= 0;
      end 
      if(_mystream_stream_oready) begin
        _mystream_sum_vec21_sink_wenable <= 0;
        _mystream_sum_vec21_sink_fifo_enq <= 0;
      end 
      if(_mystream_stream_oready) begin
        _mystream_sum_vec22_sink_wenable <= 0;
        _mystream_sum_vec22_sink_fifo_enq <= 0;
      end 
      if(_mystream_stream_oready) begin
        _mystream_sum_vec23_sink_wenable <= 0;
        _mystream_sum_vec23_sink_fifo_enq <= 0;
      end 
      if(_mystream_stream_oready) begin
        _mystream_sum_vec24_sink_wenable <= 0;
        _mystream_sum_vec24_sink_fifo_enq <= 0;
      end 
      if(_mystream_stream_oready) begin
        _mystream_sum_vec25_sink_wenable <= 0;
        _mystream_sum_vec25_sink_fifo_enq <= 0;
      end 
      if(_mystream_stream_oready) begin
        _mystream_sum_vec26_sink_wenable <= 0;
        _mystream_sum_vec26_sink_fifo_enq <= 0;
      end 
      if(_mystream_stream_oready) begin
        _mystream_sum_vec27_sink_wenable <= 0;
        _mystream_sum_vec27_sink_fifo_enq <= 0;
      end 
      if(_mystream_stream_oready) begin
        _mystream_sum_vec28_sink_wenable <= 0;
        _mystream_sum_vec28_sink_fifo_enq <= 0;
      end 
      if(_mystream_stream_oready) begin
        _mystream_sum_vec29_sink_wenable <= 0;
        _mystream_sum_vec29_sink_fifo_enq <= 0;
      end 
      if(_mystream_stream_oready) begin
        _mystream_sum_vec30_sink_wenable <= 0;
        _mystream_sum_vec30_sink_fifo_enq <= 0;
      end 
      if(_mystream_stream_oready) begin
        _mystream_sum_vec31_sink_wenable <= 0;
        _mystream_sum_vec31_sink_fifo_enq <= 0;
      end 
      if(_mystream_stream_oready) begin
        __mystream_stream_ivalid_1 <= _mystream_stream_ivalid;
      end 
      if(_mystream_stream_oready) begin
        __mystream_stream_ivalid_2 <= __mystream_stream_ivalid_1;
      end 
      if(_mystream_stream_oready) begin
        __mystream_stream_ivalid_3 <= __mystream_stream_ivalid_2;
      end 
      if(_mystream_stream_oready) begin
        __mystream_stream_ivalid_4 <= __mystream_stream_ivalid_3;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_98 <= mystream_a0_data + mystream_b0_data;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_99 <= mystream_a1_data + mystream_b1_data;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_100 <= mystream_a2_data + mystream_b2_data;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_101 <= mystream_a3_data + mystream_b3_data;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_102 <= mystream_a4_data + mystream_b4_data;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_103 <= mystream_a5_data + mystream_b5_data;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_104 <= mystream_a6_data + mystream_b6_data;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_105 <= mystream_a7_data + mystream_b7_data;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_106 <= mystream_a8_data + mystream_b8_data;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_107 <= mystream_a9_data + mystream_b9_data;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_108 <= mystream_a10_data + mystream_b10_data;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_109 <= mystream_a11_data + mystream_b11_data;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_110 <= mystream_a12_data + mystream_b12_data;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_111 <= mystream_a13_data + mystream_b13_data;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_112 <= mystream_a14_data + mystream_b14_data;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_113 <= mystream_a15_data + mystream_b15_data;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_114 <= mystream_a16_data + mystream_b16_data;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_115 <= mystream_a17_data + mystream_b17_data;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_116 <= mystream_a18_data + mystream_b18_data;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_117 <= mystream_a19_data + mystream_b19_data;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_118 <= mystream_a20_data + mystream_b20_data;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_119 <= mystream_a21_data + mystream_b21_data;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_120 <= mystream_a22_data + mystream_b22_data;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_121 <= mystream_a23_data + mystream_b23_data;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_122 <= mystream_a24_data + mystream_b24_data;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_123 <= mystream_a25_data + mystream_b25_data;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_124 <= mystream_a26_data + mystream_b26_data;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_125 <= mystream_a27_data + mystream_b27_data;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_126 <= mystream_a28_data + mystream_b28_data;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_127 <= mystream_a29_data + mystream_b29_data;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_128 <= mystream_a30_data + mystream_b30_data;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_129 <= mystream_a31_data + mystream_b31_data;
      end 
      if(_mystream_stream_ivalid && _mystream_stream_oready && _counter_reset_cond_131) begin
        _counter_data_131 <= 1'sd0;
      end 
      if(_mystream_stream_ivalid && _mystream_stream_oready) begin
        _counter_data_131 <= _counter_current_count_131;
      end 
      if(_mystream_stream_ivalid && _mystream_stream_oready) begin
        _counter_count_131 <= _counter_current_count_131 + 7'sd32;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_294__variable_1 <= mystream_tensor_size_data;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_134 <= _counter_data_131 + 1'sd0;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_137 <= _counter_data_131 + 2'sd1;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_140 <= _counter_data_131 + 3'sd2;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_143 <= _counter_data_131 + 3'sd3;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_146 <= _counter_data_131 + 4'sd4;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_149 <= _counter_data_131 + 4'sd5;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_152 <= _counter_data_131 + 4'sd6;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_155 <= _counter_data_131 + 4'sd7;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_158 <= _counter_data_131 + 5'sd8;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_161 <= _counter_data_131 + 5'sd9;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_164 <= _counter_data_131 + 5'sd10;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_167 <= _counter_data_131 + 5'sd11;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_170 <= _counter_data_131 + 5'sd12;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_173 <= _counter_data_131 + 5'sd13;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_176 <= _counter_data_131 + 5'sd14;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_179 <= _counter_data_131 + 5'sd15;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_182 <= _counter_data_131 + 6'sd16;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_185 <= _counter_data_131 + 6'sd17;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_188 <= _counter_data_131 + 6'sd18;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_191 <= _counter_data_131 + 6'sd19;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_194 <= _counter_data_131 + 6'sd20;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_197 <= _counter_data_131 + 6'sd21;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_200 <= _counter_data_131 + 6'sd22;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_203 <= _counter_data_131 + 6'sd23;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_206 <= _counter_data_131 + 6'sd24;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_209 <= _counter_data_131 + 6'sd25;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_212 <= _counter_data_131 + 6'sd26;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_215 <= _counter_data_131 + 6'sd27;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_218 <= _counter_data_131 + 6'sd28;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_221 <= _counter_data_131 + 6'sd29;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_224 <= _counter_data_131 + 6'sd30;
      end 
      if(_mystream_stream_oready) begin
        _plus_data_227 <= _counter_data_131 + 6'sd31;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_295__delay_294__variable_1 <= __delay_data_294__variable_1;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_296_plus_98 <= _plus_data_98;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_298_plus_99 <= _plus_data_99;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_300_plus_100 <= _plus_data_100;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_302_plus_101 <= _plus_data_101;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_304_plus_102 <= _plus_data_102;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_306_plus_103 <= _plus_data_103;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_308_plus_104 <= _plus_data_104;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_310_plus_105 <= _plus_data_105;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_312_plus_106 <= _plus_data_106;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_314_plus_107 <= _plus_data_107;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_316_plus_108 <= _plus_data_108;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_318_plus_109 <= _plus_data_109;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_320_plus_110 <= _plus_data_110;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_322_plus_111 <= _plus_data_111;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_324_plus_112 <= _plus_data_112;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_326_plus_113 <= _plus_data_113;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_328_plus_114 <= _plus_data_114;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_330_plus_115 <= _plus_data_115;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_332_plus_116 <= _plus_data_116;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_334_plus_117 <= _plus_data_117;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_336_plus_118 <= _plus_data_118;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_338_plus_119 <= _plus_data_119;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_340_plus_120 <= _plus_data_120;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_342_plus_121 <= _plus_data_121;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_344_plus_122 <= _plus_data_122;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_346_plus_123 <= _plus_data_123;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_348_plus_124 <= _plus_data_124;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_350_plus_125 <= _plus_data_125;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_352_plus_126 <= _plus_data_126;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_354_plus_127 <= _plus_data_127;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_356_plus_128 <= _plus_data_128;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_358_plus_129 <= _plus_data_129;
      end 
      if(_mystream_stream_oready) begin
        _greatereq_data_136 <= _plus_data_134 >= __delay_data_295__delay_294__variable_1;
      end 
      if(_mystream_stream_oready) begin
        _greatereq_data_139 <= _plus_data_137 >= __delay_data_295__delay_294__variable_1;
      end 
      if(_mystream_stream_oready) begin
        _greatereq_data_142 <= _plus_data_140 >= __delay_data_295__delay_294__variable_1;
      end 
      if(_mystream_stream_oready) begin
        _greatereq_data_145 <= _plus_data_143 >= __delay_data_295__delay_294__variable_1;
      end 
      if(_mystream_stream_oready) begin
        _greatereq_data_148 <= _plus_data_146 >= __delay_data_295__delay_294__variable_1;
      end 
      if(_mystream_stream_oready) begin
        _greatereq_data_151 <= _plus_data_149 >= __delay_data_295__delay_294__variable_1;
      end 
      if(_mystream_stream_oready) begin
        _greatereq_data_154 <= _plus_data_152 >= __delay_data_295__delay_294__variable_1;
      end 
      if(_mystream_stream_oready) begin
        _greatereq_data_157 <= _plus_data_155 >= __delay_data_295__delay_294__variable_1;
      end 
      if(_mystream_stream_oready) begin
        _greatereq_data_160 <= _plus_data_158 >= __delay_data_295__delay_294__variable_1;
      end 
      if(_mystream_stream_oready) begin
        _greatereq_data_163 <= _plus_data_161 >= __delay_data_295__delay_294__variable_1;
      end 
      if(_mystream_stream_oready) begin
        _greatereq_data_166 <= _plus_data_164 >= __delay_data_295__delay_294__variable_1;
      end 
      if(_mystream_stream_oready) begin
        _greatereq_data_169 <= _plus_data_167 >= __delay_data_295__delay_294__variable_1;
      end 
      if(_mystream_stream_oready) begin
        _greatereq_data_172 <= _plus_data_170 >= __delay_data_295__delay_294__variable_1;
      end 
      if(_mystream_stream_oready) begin
        _greatereq_data_175 <= _plus_data_173 >= __delay_data_295__delay_294__variable_1;
      end 
      if(_mystream_stream_oready) begin
        _greatereq_data_178 <= _plus_data_176 >= __delay_data_295__delay_294__variable_1;
      end 
      if(_mystream_stream_oready) begin
        _greatereq_data_181 <= _plus_data_179 >= __delay_data_295__delay_294__variable_1;
      end 
      if(_mystream_stream_oready) begin
        _greatereq_data_184 <= _plus_data_182 >= __delay_data_295__delay_294__variable_1;
      end 
      if(_mystream_stream_oready) begin
        _greatereq_data_187 <= _plus_data_185 >= __delay_data_295__delay_294__variable_1;
      end 
      if(_mystream_stream_oready) begin
        _greatereq_data_190 <= _plus_data_188 >= __delay_data_295__delay_294__variable_1;
      end 
      if(_mystream_stream_oready) begin
        _greatereq_data_193 <= _plus_data_191 >= __delay_data_295__delay_294__variable_1;
      end 
      if(_mystream_stream_oready) begin
        _greatereq_data_196 <= _plus_data_194 >= __delay_data_295__delay_294__variable_1;
      end 
      if(_mystream_stream_oready) begin
        _greatereq_data_199 <= _plus_data_197 >= __delay_data_295__delay_294__variable_1;
      end 
      if(_mystream_stream_oready) begin
        _greatereq_data_202 <= _plus_data_200 >= __delay_data_295__delay_294__variable_1;
      end 
      if(_mystream_stream_oready) begin
        _greatereq_data_205 <= _plus_data_203 >= __delay_data_295__delay_294__variable_1;
      end 
      if(_mystream_stream_oready) begin
        _greatereq_data_208 <= _plus_data_206 >= __delay_data_295__delay_294__variable_1;
      end 
      if(_mystream_stream_oready) begin
        _greatereq_data_211 <= _plus_data_209 >= __delay_data_295__delay_294__variable_1;
      end 
      if(_mystream_stream_oready) begin
        _greatereq_data_214 <= _plus_data_212 >= __delay_data_295__delay_294__variable_1;
      end 
      if(_mystream_stream_oready) begin
        _greatereq_data_217 <= _plus_data_215 >= __delay_data_295__delay_294__variable_1;
      end 
      if(_mystream_stream_oready) begin
        _greatereq_data_220 <= _plus_data_218 >= __delay_data_295__delay_294__variable_1;
      end 
      if(_mystream_stream_oready) begin
        _greatereq_data_223 <= _plus_data_221 >= __delay_data_295__delay_294__variable_1;
      end 
      if(_mystream_stream_oready) begin
        _greatereq_data_226 <= _plus_data_224 >= __delay_data_295__delay_294__variable_1;
      end 
      if(_mystream_stream_oready) begin
        _greatereq_data_229 <= _plus_data_227 >= __delay_data_295__delay_294__variable_1;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_297__delay_296_plus_98 <= __delay_data_296_plus_98;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_299__delay_298_plus_99 <= __delay_data_298_plus_99;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_301__delay_300_plus_100 <= __delay_data_300_plus_100;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_303__delay_302_plus_101 <= __delay_data_302_plus_101;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_305__delay_304_plus_102 <= __delay_data_304_plus_102;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_307__delay_306_plus_103 <= __delay_data_306_plus_103;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_309__delay_308_plus_104 <= __delay_data_308_plus_104;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_311__delay_310_plus_105 <= __delay_data_310_plus_105;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_313__delay_312_plus_106 <= __delay_data_312_plus_106;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_315__delay_314_plus_107 <= __delay_data_314_plus_107;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_317__delay_316_plus_108 <= __delay_data_316_plus_108;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_319__delay_318_plus_109 <= __delay_data_318_plus_109;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_321__delay_320_plus_110 <= __delay_data_320_plus_110;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_323__delay_322_plus_111 <= __delay_data_322_plus_111;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_325__delay_324_plus_112 <= __delay_data_324_plus_112;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_327__delay_326_plus_113 <= __delay_data_326_plus_113;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_329__delay_328_plus_114 <= __delay_data_328_plus_114;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_331__delay_330_plus_115 <= __delay_data_330_plus_115;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_333__delay_332_plus_116 <= __delay_data_332_plus_116;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_335__delay_334_plus_117 <= __delay_data_334_plus_117;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_337__delay_336_plus_118 <= __delay_data_336_plus_118;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_339__delay_338_plus_119 <= __delay_data_338_plus_119;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_341__delay_340_plus_120 <= __delay_data_340_plus_120;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_343__delay_342_plus_121 <= __delay_data_342_plus_121;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_345__delay_344_plus_122 <= __delay_data_344_plus_122;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_347__delay_346_plus_123 <= __delay_data_346_plus_123;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_349__delay_348_plus_124 <= __delay_data_348_plus_124;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_351__delay_350_plus_125 <= __delay_data_350_plus_125;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_353__delay_352_plus_126 <= __delay_data_352_plus_126;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_355__delay_354_plus_127 <= __delay_data_354_plus_127;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_357__delay_356_plus_128 <= __delay_data_356_plus_128;
      end 
      if(_mystream_stream_oready) begin
        __delay_data_359__delay_358_plus_129 <= __delay_data_358_plus_129;
      end 
      if(_mystream_stream_oready) begin
        _cond_data_230 <= (_greatereq_data_136)? 1'sd0 : __delay_data_297__delay_296_plus_98;
      end 
      if(_mystream_stream_oready) begin
        _cond_data_232 <= (_greatereq_data_139)? 1'sd0 : __delay_data_299__delay_298_plus_99;
      end 
      if(_mystream_stream_oready) begin
        _cond_data_234 <= (_greatereq_data_142)? 1'sd0 : __delay_data_301__delay_300_plus_100;
      end 
      if(_mystream_stream_oready) begin
        _cond_data_236 <= (_greatereq_data_145)? 1'sd0 : __delay_data_303__delay_302_plus_101;
      end 
      if(_mystream_stream_oready) begin
        _cond_data_238 <= (_greatereq_data_148)? 1'sd0 : __delay_data_305__delay_304_plus_102;
      end 
      if(_mystream_stream_oready) begin
        _cond_data_240 <= (_greatereq_data_151)? 1'sd0 : __delay_data_307__delay_306_plus_103;
      end 
      if(_mystream_stream_oready) begin
        _cond_data_242 <= (_greatereq_data_154)? 1'sd0 : __delay_data_309__delay_308_plus_104;
      end 
      if(_mystream_stream_oready) begin
        _cond_data_244 <= (_greatereq_data_157)? 1'sd0 : __delay_data_311__delay_310_plus_105;
      end 
      if(_mystream_stream_oready) begin
        _cond_data_246 <= (_greatereq_data_160)? 1'sd0 : __delay_data_313__delay_312_plus_106;
      end 
      if(_mystream_stream_oready) begin
        _cond_data_248 <= (_greatereq_data_163)? 1'sd0 : __delay_data_315__delay_314_plus_107;
      end 
      if(_mystream_stream_oready) begin
        _cond_data_250 <= (_greatereq_data_166)? 1'sd0 : __delay_data_317__delay_316_plus_108;
      end 
      if(_mystream_stream_oready) begin
        _cond_data_252 <= (_greatereq_data_169)? 1'sd0 : __delay_data_319__delay_318_plus_109;
      end 
      if(_mystream_stream_oready) begin
        _cond_data_254 <= (_greatereq_data_172)? 1'sd0 : __delay_data_321__delay_320_plus_110;
      end 
      if(_mystream_stream_oready) begin
        _cond_data_256 <= (_greatereq_data_175)? 1'sd0 : __delay_data_323__delay_322_plus_111;
      end 
      if(_mystream_stream_oready) begin
        _cond_data_258 <= (_greatereq_data_178)? 1'sd0 : __delay_data_325__delay_324_plus_112;
      end 
      if(_mystream_stream_oready) begin
        _cond_data_260 <= (_greatereq_data_181)? 1'sd0 : __delay_data_327__delay_326_plus_113;
      end 
      if(_mystream_stream_oready) begin
        _cond_data_262 <= (_greatereq_data_184)? 1'sd0 : __delay_data_329__delay_328_plus_114;
      end 
      if(_mystream_stream_oready) begin
        _cond_data_264 <= (_greatereq_data_187)? 1'sd0 : __delay_data_331__delay_330_plus_115;
      end 
      if(_mystream_stream_oready) begin
        _cond_data_266 <= (_greatereq_data_190)? 1'sd0 : __delay_data_333__delay_332_plus_116;
      end 
      if(_mystream_stream_oready) begin
        _cond_data_268 <= (_greatereq_data_193)? 1'sd0 : __delay_data_335__delay_334_plus_117;
      end 
      if(_mystream_stream_oready) begin
        _cond_data_270 <= (_greatereq_data_196)? 1'sd0 : __delay_data_337__delay_336_plus_118;
      end 
      if(_mystream_stream_oready) begin
        _cond_data_272 <= (_greatereq_data_199)? 1'sd0 : __delay_data_339__delay_338_plus_119;
      end 
      if(_mystream_stream_oready) begin
        _cond_data_274 <= (_greatereq_data_202)? 1'sd0 : __delay_data_341__delay_340_plus_120;
      end 
      if(_mystream_stream_oready) begin
        _cond_data_276 <= (_greatereq_data_205)? 1'sd0 : __delay_data_343__delay_342_plus_121;
      end 
      if(_mystream_stream_oready) begin
        _cond_data_278 <= (_greatereq_data_208)? 1'sd0 : __delay_data_345__delay_344_plus_122;
      end 
      if(_mystream_stream_oready) begin
        _cond_data_280 <= (_greatereq_data_211)? 1'sd0 : __delay_data_347__delay_346_plus_123;
      end 
      if(_mystream_stream_oready) begin
        _cond_data_282 <= (_greatereq_data_214)? 1'sd0 : __delay_data_349__delay_348_plus_124;
      end 
      if(_mystream_stream_oready) begin
        _cond_data_284 <= (_greatereq_data_217)? 1'sd0 : __delay_data_351__delay_350_plus_125;
      end 
      if(_mystream_stream_oready) begin
        _cond_data_286 <= (_greatereq_data_220)? 1'sd0 : __delay_data_353__delay_352_plus_126;
      end 
      if(_mystream_stream_oready) begin
        _cond_data_288 <= (_greatereq_data_223)? 1'sd0 : __delay_data_355__delay_354_plus_127;
      end 
      if(_mystream_stream_oready) begin
        _cond_data_290 <= (_greatereq_data_226)? 1'sd0 : __delay_data_357__delay_356_plus_128;
      end 
      if(_mystream_stream_oready) begin
        _cond_data_292 <= (_greatereq_data_229)? 1'sd0 : __delay_data_359__delay_358_plus_129;
      end 
      if(_set_flag_183) begin
        _mystream_tensor_size_next_parameter_data <= _th_comp_size_3;
      end 
      if(_mystream_source_start) begin
        __variable_wdata_1 <= _mystream_tensor_size_next_parameter_data;
      end 
      if(_set_flag_184) begin
        _mystream_size_next_parameter_data <= _th_comp_size_3 + 32 - 1 >>> 5;
      end 
      if(_mystream_source_start) begin
        __variable_wdata_0 <= _mystream_size_next_parameter_data;
      end 
      if(_set_flag_185) begin
        _mystream_a0_source_mode <= 5'b1;
        _mystream_a0_source_offset <= _th_comp_offset_4;
        _mystream_a0_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_a0_source_stride <= 1;
      end 
      if(_set_flag_185) begin
        _mystream_a0_source_sel <= 1;
      end 
      if(_mystream_source_start && _mystream_a0_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_a0_source_offset_buf <= _mystream_a0_source_offset;
        _mystream_a0_source_size_buf <= _mystream_a0_source_size;
        _mystream_a0_source_stride_buf <= _mystream_a0_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_2 <= _mystream_a0_source_ram_rdata;
      end 
      if((_mystream_a0_source_fsm_0 == 1) && _mystream_stream_oready) begin
        _mystream_a0_idle <= 0;
        _mystream_a0_source_ram_raddr <= _mystream_a0_source_offset_buf;
        _mystream_a0_source_ram_renable <= 1;
        _mystream_a0_source_count <= _mystream_a0_source_size_buf;
      end 
      if((_mystream_a0_source_fsm_0 == 2) && _mystream_stream_oready) begin
        _mystream_a0_source_ram_raddr <= _mystream_a0_source_ram_raddr + _mystream_a0_source_stride_buf;
        _mystream_a0_source_ram_renable <= 1;
        _mystream_a0_source_count <= _mystream_a0_source_count - 1;
      end 
      if((_mystream_a0_source_fsm_0 == 2) && (_mystream_a0_source_count == 1) && _mystream_stream_oready) begin
        _mystream_a0_source_ram_renable <= 0;
        _mystream_a0_idle <= 1;
      end 
      if((_mystream_a0_source_fsm_0 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_a0_source_ram_renable <= 0;
        _mystream_a0_idle <= 1;
      end 
      if(_set_flag_188) begin
        _mystream_a1_source_mode <= 5'b1;
        _mystream_a1_source_offset <= _th_comp_offset_4;
        _mystream_a1_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_a1_source_stride <= 1;
      end 
      if(_set_flag_188) begin
        _mystream_a1_source_sel <= 2;
      end 
      if(_mystream_source_start && _mystream_a1_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_a1_source_offset_buf <= _mystream_a1_source_offset;
        _mystream_a1_source_size_buf <= _mystream_a1_source_size;
        _mystream_a1_source_stride_buf <= _mystream_a1_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_3 <= _mystream_a1_source_ram_rdata;
      end 
      if((_mystream_a1_source_fsm_1 == 1) && _mystream_stream_oready) begin
        _mystream_a1_idle <= 0;
        _mystream_a1_source_ram_raddr <= _mystream_a1_source_offset_buf;
        _mystream_a1_source_ram_renable <= 1;
        _mystream_a1_source_count <= _mystream_a1_source_size_buf;
      end 
      if((_mystream_a1_source_fsm_1 == 2) && _mystream_stream_oready) begin
        _mystream_a1_source_ram_raddr <= _mystream_a1_source_ram_raddr + _mystream_a1_source_stride_buf;
        _mystream_a1_source_ram_renable <= 1;
        _mystream_a1_source_count <= _mystream_a1_source_count - 1;
      end 
      if((_mystream_a1_source_fsm_1 == 2) && (_mystream_a1_source_count == 1) && _mystream_stream_oready) begin
        _mystream_a1_source_ram_renable <= 0;
        _mystream_a1_idle <= 1;
      end 
      if((_mystream_a1_source_fsm_1 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_a1_source_ram_renable <= 0;
        _mystream_a1_idle <= 1;
      end 
      if(_set_flag_191) begin
        _mystream_a2_source_mode <= 5'b1;
        _mystream_a2_source_offset <= _th_comp_offset_4;
        _mystream_a2_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_a2_source_stride <= 1;
      end 
      if(_set_flag_191) begin
        _mystream_a2_source_sel <= 3;
      end 
      if(_mystream_source_start && _mystream_a2_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_a2_source_offset_buf <= _mystream_a2_source_offset;
        _mystream_a2_source_size_buf <= _mystream_a2_source_size;
        _mystream_a2_source_stride_buf <= _mystream_a2_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_4 <= _mystream_a2_source_ram_rdata;
      end 
      if((_mystream_a2_source_fsm_2 == 1) && _mystream_stream_oready) begin
        _mystream_a2_idle <= 0;
        _mystream_a2_source_ram_raddr <= _mystream_a2_source_offset_buf;
        _mystream_a2_source_ram_renable <= 1;
        _mystream_a2_source_count <= _mystream_a2_source_size_buf;
      end 
      if((_mystream_a2_source_fsm_2 == 2) && _mystream_stream_oready) begin
        _mystream_a2_source_ram_raddr <= _mystream_a2_source_ram_raddr + _mystream_a2_source_stride_buf;
        _mystream_a2_source_ram_renable <= 1;
        _mystream_a2_source_count <= _mystream_a2_source_count - 1;
      end 
      if((_mystream_a2_source_fsm_2 == 2) && (_mystream_a2_source_count == 1) && _mystream_stream_oready) begin
        _mystream_a2_source_ram_renable <= 0;
        _mystream_a2_idle <= 1;
      end 
      if((_mystream_a2_source_fsm_2 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_a2_source_ram_renable <= 0;
        _mystream_a2_idle <= 1;
      end 
      if(_set_flag_194) begin
        _mystream_a3_source_mode <= 5'b1;
        _mystream_a3_source_offset <= _th_comp_offset_4;
        _mystream_a3_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_a3_source_stride <= 1;
      end 
      if(_set_flag_194) begin
        _mystream_a3_source_sel <= 4;
      end 
      if(_mystream_source_start && _mystream_a3_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_a3_source_offset_buf <= _mystream_a3_source_offset;
        _mystream_a3_source_size_buf <= _mystream_a3_source_size;
        _mystream_a3_source_stride_buf <= _mystream_a3_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_5 <= _mystream_a3_source_ram_rdata;
      end 
      if((_mystream_a3_source_fsm_3 == 1) && _mystream_stream_oready) begin
        _mystream_a3_idle <= 0;
        _mystream_a3_source_ram_raddr <= _mystream_a3_source_offset_buf;
        _mystream_a3_source_ram_renable <= 1;
        _mystream_a3_source_count <= _mystream_a3_source_size_buf;
      end 
      if((_mystream_a3_source_fsm_3 == 2) && _mystream_stream_oready) begin
        _mystream_a3_source_ram_raddr <= _mystream_a3_source_ram_raddr + _mystream_a3_source_stride_buf;
        _mystream_a3_source_ram_renable <= 1;
        _mystream_a3_source_count <= _mystream_a3_source_count - 1;
      end 
      if((_mystream_a3_source_fsm_3 == 2) && (_mystream_a3_source_count == 1) && _mystream_stream_oready) begin
        _mystream_a3_source_ram_renable <= 0;
        _mystream_a3_idle <= 1;
      end 
      if((_mystream_a3_source_fsm_3 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_a3_source_ram_renable <= 0;
        _mystream_a3_idle <= 1;
      end 
      if(_set_flag_197) begin
        _mystream_a4_source_mode <= 5'b1;
        _mystream_a4_source_offset <= _th_comp_offset_4;
        _mystream_a4_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_a4_source_stride <= 1;
      end 
      if(_set_flag_197) begin
        _mystream_a4_source_sel <= 5;
      end 
      if(_mystream_source_start && _mystream_a4_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_a4_source_offset_buf <= _mystream_a4_source_offset;
        _mystream_a4_source_size_buf <= _mystream_a4_source_size;
        _mystream_a4_source_stride_buf <= _mystream_a4_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_6 <= _mystream_a4_source_ram_rdata;
      end 
      if((_mystream_a4_source_fsm_4 == 1) && _mystream_stream_oready) begin
        _mystream_a4_idle <= 0;
        _mystream_a4_source_ram_raddr <= _mystream_a4_source_offset_buf;
        _mystream_a4_source_ram_renable <= 1;
        _mystream_a4_source_count <= _mystream_a4_source_size_buf;
      end 
      if((_mystream_a4_source_fsm_4 == 2) && _mystream_stream_oready) begin
        _mystream_a4_source_ram_raddr <= _mystream_a4_source_ram_raddr + _mystream_a4_source_stride_buf;
        _mystream_a4_source_ram_renable <= 1;
        _mystream_a4_source_count <= _mystream_a4_source_count - 1;
      end 
      if((_mystream_a4_source_fsm_4 == 2) && (_mystream_a4_source_count == 1) && _mystream_stream_oready) begin
        _mystream_a4_source_ram_renable <= 0;
        _mystream_a4_idle <= 1;
      end 
      if((_mystream_a4_source_fsm_4 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_a4_source_ram_renable <= 0;
        _mystream_a4_idle <= 1;
      end 
      if(_set_flag_200) begin
        _mystream_a5_source_mode <= 5'b1;
        _mystream_a5_source_offset <= _th_comp_offset_4;
        _mystream_a5_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_a5_source_stride <= 1;
      end 
      if(_set_flag_200) begin
        _mystream_a5_source_sel <= 6;
      end 
      if(_mystream_source_start && _mystream_a5_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_a5_source_offset_buf <= _mystream_a5_source_offset;
        _mystream_a5_source_size_buf <= _mystream_a5_source_size;
        _mystream_a5_source_stride_buf <= _mystream_a5_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_7 <= _mystream_a5_source_ram_rdata;
      end 
      if((_mystream_a5_source_fsm_5 == 1) && _mystream_stream_oready) begin
        _mystream_a5_idle <= 0;
        _mystream_a5_source_ram_raddr <= _mystream_a5_source_offset_buf;
        _mystream_a5_source_ram_renable <= 1;
        _mystream_a5_source_count <= _mystream_a5_source_size_buf;
      end 
      if((_mystream_a5_source_fsm_5 == 2) && _mystream_stream_oready) begin
        _mystream_a5_source_ram_raddr <= _mystream_a5_source_ram_raddr + _mystream_a5_source_stride_buf;
        _mystream_a5_source_ram_renable <= 1;
        _mystream_a5_source_count <= _mystream_a5_source_count - 1;
      end 
      if((_mystream_a5_source_fsm_5 == 2) && (_mystream_a5_source_count == 1) && _mystream_stream_oready) begin
        _mystream_a5_source_ram_renable <= 0;
        _mystream_a5_idle <= 1;
      end 
      if((_mystream_a5_source_fsm_5 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_a5_source_ram_renable <= 0;
        _mystream_a5_idle <= 1;
      end 
      if(_set_flag_203) begin
        _mystream_a6_source_mode <= 5'b1;
        _mystream_a6_source_offset <= _th_comp_offset_4;
        _mystream_a6_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_a6_source_stride <= 1;
      end 
      if(_set_flag_203) begin
        _mystream_a6_source_sel <= 7;
      end 
      if(_mystream_source_start && _mystream_a6_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_a6_source_offset_buf <= _mystream_a6_source_offset;
        _mystream_a6_source_size_buf <= _mystream_a6_source_size;
        _mystream_a6_source_stride_buf <= _mystream_a6_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_8 <= _mystream_a6_source_ram_rdata;
      end 
      if((_mystream_a6_source_fsm_6 == 1) && _mystream_stream_oready) begin
        _mystream_a6_idle <= 0;
        _mystream_a6_source_ram_raddr <= _mystream_a6_source_offset_buf;
        _mystream_a6_source_ram_renable <= 1;
        _mystream_a6_source_count <= _mystream_a6_source_size_buf;
      end 
      if((_mystream_a6_source_fsm_6 == 2) && _mystream_stream_oready) begin
        _mystream_a6_source_ram_raddr <= _mystream_a6_source_ram_raddr + _mystream_a6_source_stride_buf;
        _mystream_a6_source_ram_renable <= 1;
        _mystream_a6_source_count <= _mystream_a6_source_count - 1;
      end 
      if((_mystream_a6_source_fsm_6 == 2) && (_mystream_a6_source_count == 1) && _mystream_stream_oready) begin
        _mystream_a6_source_ram_renable <= 0;
        _mystream_a6_idle <= 1;
      end 
      if((_mystream_a6_source_fsm_6 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_a6_source_ram_renable <= 0;
        _mystream_a6_idle <= 1;
      end 
      if(_set_flag_206) begin
        _mystream_a7_source_mode <= 5'b1;
        _mystream_a7_source_offset <= _th_comp_offset_4;
        _mystream_a7_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_a7_source_stride <= 1;
      end 
      if(_set_flag_206) begin
        _mystream_a7_source_sel <= 8;
      end 
      if(_mystream_source_start && _mystream_a7_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_a7_source_offset_buf <= _mystream_a7_source_offset;
        _mystream_a7_source_size_buf <= _mystream_a7_source_size;
        _mystream_a7_source_stride_buf <= _mystream_a7_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_9 <= _mystream_a7_source_ram_rdata;
      end 
      if((_mystream_a7_source_fsm_7 == 1) && _mystream_stream_oready) begin
        _mystream_a7_idle <= 0;
        _mystream_a7_source_ram_raddr <= _mystream_a7_source_offset_buf;
        _mystream_a7_source_ram_renable <= 1;
        _mystream_a7_source_count <= _mystream_a7_source_size_buf;
      end 
      if((_mystream_a7_source_fsm_7 == 2) && _mystream_stream_oready) begin
        _mystream_a7_source_ram_raddr <= _mystream_a7_source_ram_raddr + _mystream_a7_source_stride_buf;
        _mystream_a7_source_ram_renable <= 1;
        _mystream_a7_source_count <= _mystream_a7_source_count - 1;
      end 
      if((_mystream_a7_source_fsm_7 == 2) && (_mystream_a7_source_count == 1) && _mystream_stream_oready) begin
        _mystream_a7_source_ram_renable <= 0;
        _mystream_a7_idle <= 1;
      end 
      if((_mystream_a7_source_fsm_7 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_a7_source_ram_renable <= 0;
        _mystream_a7_idle <= 1;
      end 
      if(_set_flag_209) begin
        _mystream_a8_source_mode <= 5'b1;
        _mystream_a8_source_offset <= _th_comp_offset_4;
        _mystream_a8_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_a8_source_stride <= 1;
      end 
      if(_set_flag_209) begin
        _mystream_a8_source_sel <= 9;
      end 
      if(_mystream_source_start && _mystream_a8_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_a8_source_offset_buf <= _mystream_a8_source_offset;
        _mystream_a8_source_size_buf <= _mystream_a8_source_size;
        _mystream_a8_source_stride_buf <= _mystream_a8_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_10 <= _mystream_a8_source_ram_rdata;
      end 
      if((_mystream_a8_source_fsm_8 == 1) && _mystream_stream_oready) begin
        _mystream_a8_idle <= 0;
        _mystream_a8_source_ram_raddr <= _mystream_a8_source_offset_buf;
        _mystream_a8_source_ram_renable <= 1;
        _mystream_a8_source_count <= _mystream_a8_source_size_buf;
      end 
      if((_mystream_a8_source_fsm_8 == 2) && _mystream_stream_oready) begin
        _mystream_a8_source_ram_raddr <= _mystream_a8_source_ram_raddr + _mystream_a8_source_stride_buf;
        _mystream_a8_source_ram_renable <= 1;
        _mystream_a8_source_count <= _mystream_a8_source_count - 1;
      end 
      if((_mystream_a8_source_fsm_8 == 2) && (_mystream_a8_source_count == 1) && _mystream_stream_oready) begin
        _mystream_a8_source_ram_renable <= 0;
        _mystream_a8_idle <= 1;
      end 
      if((_mystream_a8_source_fsm_8 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_a8_source_ram_renable <= 0;
        _mystream_a8_idle <= 1;
      end 
      if(_set_flag_212) begin
        _mystream_a9_source_mode <= 5'b1;
        _mystream_a9_source_offset <= _th_comp_offset_4;
        _mystream_a9_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_a9_source_stride <= 1;
      end 
      if(_set_flag_212) begin
        _mystream_a9_source_sel <= 10;
      end 
      if(_mystream_source_start && _mystream_a9_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_a9_source_offset_buf <= _mystream_a9_source_offset;
        _mystream_a9_source_size_buf <= _mystream_a9_source_size;
        _mystream_a9_source_stride_buf <= _mystream_a9_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_11 <= _mystream_a9_source_ram_rdata;
      end 
      if((_mystream_a9_source_fsm_9 == 1) && _mystream_stream_oready) begin
        _mystream_a9_idle <= 0;
        _mystream_a9_source_ram_raddr <= _mystream_a9_source_offset_buf;
        _mystream_a9_source_ram_renable <= 1;
        _mystream_a9_source_count <= _mystream_a9_source_size_buf;
      end 
      if((_mystream_a9_source_fsm_9 == 2) && _mystream_stream_oready) begin
        _mystream_a9_source_ram_raddr <= _mystream_a9_source_ram_raddr + _mystream_a9_source_stride_buf;
        _mystream_a9_source_ram_renable <= 1;
        _mystream_a9_source_count <= _mystream_a9_source_count - 1;
      end 
      if((_mystream_a9_source_fsm_9 == 2) && (_mystream_a9_source_count == 1) && _mystream_stream_oready) begin
        _mystream_a9_source_ram_renable <= 0;
        _mystream_a9_idle <= 1;
      end 
      if((_mystream_a9_source_fsm_9 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_a9_source_ram_renable <= 0;
        _mystream_a9_idle <= 1;
      end 
      if(_set_flag_215) begin
        _mystream_a10_source_mode <= 5'b1;
        _mystream_a10_source_offset <= _th_comp_offset_4;
        _mystream_a10_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_a10_source_stride <= 1;
      end 
      if(_set_flag_215) begin
        _mystream_a10_source_sel <= 11;
      end 
      if(_mystream_source_start && _mystream_a10_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_a10_source_offset_buf <= _mystream_a10_source_offset;
        _mystream_a10_source_size_buf <= _mystream_a10_source_size;
        _mystream_a10_source_stride_buf <= _mystream_a10_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_12 <= _mystream_a10_source_ram_rdata;
      end 
      if((_mystream_a10_source_fsm_10 == 1) && _mystream_stream_oready) begin
        _mystream_a10_idle <= 0;
        _mystream_a10_source_ram_raddr <= _mystream_a10_source_offset_buf;
        _mystream_a10_source_ram_renable <= 1;
        _mystream_a10_source_count <= _mystream_a10_source_size_buf;
      end 
      if((_mystream_a10_source_fsm_10 == 2) && _mystream_stream_oready) begin
        _mystream_a10_source_ram_raddr <= _mystream_a10_source_ram_raddr + _mystream_a10_source_stride_buf;
        _mystream_a10_source_ram_renable <= 1;
        _mystream_a10_source_count <= _mystream_a10_source_count - 1;
      end 
      if((_mystream_a10_source_fsm_10 == 2) && (_mystream_a10_source_count == 1) && _mystream_stream_oready) begin
        _mystream_a10_source_ram_renable <= 0;
        _mystream_a10_idle <= 1;
      end 
      if((_mystream_a10_source_fsm_10 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_a10_source_ram_renable <= 0;
        _mystream_a10_idle <= 1;
      end 
      if(_set_flag_218) begin
        _mystream_a11_source_mode <= 5'b1;
        _mystream_a11_source_offset <= _th_comp_offset_4;
        _mystream_a11_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_a11_source_stride <= 1;
      end 
      if(_set_flag_218) begin
        _mystream_a11_source_sel <= 12;
      end 
      if(_mystream_source_start && _mystream_a11_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_a11_source_offset_buf <= _mystream_a11_source_offset;
        _mystream_a11_source_size_buf <= _mystream_a11_source_size;
        _mystream_a11_source_stride_buf <= _mystream_a11_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_13 <= _mystream_a11_source_ram_rdata;
      end 
      if((_mystream_a11_source_fsm_11 == 1) && _mystream_stream_oready) begin
        _mystream_a11_idle <= 0;
        _mystream_a11_source_ram_raddr <= _mystream_a11_source_offset_buf;
        _mystream_a11_source_ram_renable <= 1;
        _mystream_a11_source_count <= _mystream_a11_source_size_buf;
      end 
      if((_mystream_a11_source_fsm_11 == 2) && _mystream_stream_oready) begin
        _mystream_a11_source_ram_raddr <= _mystream_a11_source_ram_raddr + _mystream_a11_source_stride_buf;
        _mystream_a11_source_ram_renable <= 1;
        _mystream_a11_source_count <= _mystream_a11_source_count - 1;
      end 
      if((_mystream_a11_source_fsm_11 == 2) && (_mystream_a11_source_count == 1) && _mystream_stream_oready) begin
        _mystream_a11_source_ram_renable <= 0;
        _mystream_a11_idle <= 1;
      end 
      if((_mystream_a11_source_fsm_11 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_a11_source_ram_renable <= 0;
        _mystream_a11_idle <= 1;
      end 
      if(_set_flag_221) begin
        _mystream_a12_source_mode <= 5'b1;
        _mystream_a12_source_offset <= _th_comp_offset_4;
        _mystream_a12_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_a12_source_stride <= 1;
      end 
      if(_set_flag_221) begin
        _mystream_a12_source_sel <= 13;
      end 
      if(_mystream_source_start && _mystream_a12_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_a12_source_offset_buf <= _mystream_a12_source_offset;
        _mystream_a12_source_size_buf <= _mystream_a12_source_size;
        _mystream_a12_source_stride_buf <= _mystream_a12_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_14 <= _mystream_a12_source_ram_rdata;
      end 
      if((_mystream_a12_source_fsm_12 == 1) && _mystream_stream_oready) begin
        _mystream_a12_idle <= 0;
        _mystream_a12_source_ram_raddr <= _mystream_a12_source_offset_buf;
        _mystream_a12_source_ram_renable <= 1;
        _mystream_a12_source_count <= _mystream_a12_source_size_buf;
      end 
      if((_mystream_a12_source_fsm_12 == 2) && _mystream_stream_oready) begin
        _mystream_a12_source_ram_raddr <= _mystream_a12_source_ram_raddr + _mystream_a12_source_stride_buf;
        _mystream_a12_source_ram_renable <= 1;
        _mystream_a12_source_count <= _mystream_a12_source_count - 1;
      end 
      if((_mystream_a12_source_fsm_12 == 2) && (_mystream_a12_source_count == 1) && _mystream_stream_oready) begin
        _mystream_a12_source_ram_renable <= 0;
        _mystream_a12_idle <= 1;
      end 
      if((_mystream_a12_source_fsm_12 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_a12_source_ram_renable <= 0;
        _mystream_a12_idle <= 1;
      end 
      if(_set_flag_224) begin
        _mystream_a13_source_mode <= 5'b1;
        _mystream_a13_source_offset <= _th_comp_offset_4;
        _mystream_a13_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_a13_source_stride <= 1;
      end 
      if(_set_flag_224) begin
        _mystream_a13_source_sel <= 14;
      end 
      if(_mystream_source_start && _mystream_a13_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_a13_source_offset_buf <= _mystream_a13_source_offset;
        _mystream_a13_source_size_buf <= _mystream_a13_source_size;
        _mystream_a13_source_stride_buf <= _mystream_a13_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_15 <= _mystream_a13_source_ram_rdata;
      end 
      if((_mystream_a13_source_fsm_13 == 1) && _mystream_stream_oready) begin
        _mystream_a13_idle <= 0;
        _mystream_a13_source_ram_raddr <= _mystream_a13_source_offset_buf;
        _mystream_a13_source_ram_renable <= 1;
        _mystream_a13_source_count <= _mystream_a13_source_size_buf;
      end 
      if((_mystream_a13_source_fsm_13 == 2) && _mystream_stream_oready) begin
        _mystream_a13_source_ram_raddr <= _mystream_a13_source_ram_raddr + _mystream_a13_source_stride_buf;
        _mystream_a13_source_ram_renable <= 1;
        _mystream_a13_source_count <= _mystream_a13_source_count - 1;
      end 
      if((_mystream_a13_source_fsm_13 == 2) && (_mystream_a13_source_count == 1) && _mystream_stream_oready) begin
        _mystream_a13_source_ram_renable <= 0;
        _mystream_a13_idle <= 1;
      end 
      if((_mystream_a13_source_fsm_13 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_a13_source_ram_renable <= 0;
        _mystream_a13_idle <= 1;
      end 
      if(_set_flag_227) begin
        _mystream_a14_source_mode <= 5'b1;
        _mystream_a14_source_offset <= _th_comp_offset_4;
        _mystream_a14_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_a14_source_stride <= 1;
      end 
      if(_set_flag_227) begin
        _mystream_a14_source_sel <= 15;
      end 
      if(_mystream_source_start && _mystream_a14_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_a14_source_offset_buf <= _mystream_a14_source_offset;
        _mystream_a14_source_size_buf <= _mystream_a14_source_size;
        _mystream_a14_source_stride_buf <= _mystream_a14_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_16 <= _mystream_a14_source_ram_rdata;
      end 
      if((_mystream_a14_source_fsm_14 == 1) && _mystream_stream_oready) begin
        _mystream_a14_idle <= 0;
        _mystream_a14_source_ram_raddr <= _mystream_a14_source_offset_buf;
        _mystream_a14_source_ram_renable <= 1;
        _mystream_a14_source_count <= _mystream_a14_source_size_buf;
      end 
      if((_mystream_a14_source_fsm_14 == 2) && _mystream_stream_oready) begin
        _mystream_a14_source_ram_raddr <= _mystream_a14_source_ram_raddr + _mystream_a14_source_stride_buf;
        _mystream_a14_source_ram_renable <= 1;
        _mystream_a14_source_count <= _mystream_a14_source_count - 1;
      end 
      if((_mystream_a14_source_fsm_14 == 2) && (_mystream_a14_source_count == 1) && _mystream_stream_oready) begin
        _mystream_a14_source_ram_renable <= 0;
        _mystream_a14_idle <= 1;
      end 
      if((_mystream_a14_source_fsm_14 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_a14_source_ram_renable <= 0;
        _mystream_a14_idle <= 1;
      end 
      if(_set_flag_230) begin
        _mystream_a15_source_mode <= 5'b1;
        _mystream_a15_source_offset <= _th_comp_offset_4;
        _mystream_a15_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_a15_source_stride <= 1;
      end 
      if(_set_flag_230) begin
        _mystream_a15_source_sel <= 16;
      end 
      if(_mystream_source_start && _mystream_a15_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_a15_source_offset_buf <= _mystream_a15_source_offset;
        _mystream_a15_source_size_buf <= _mystream_a15_source_size;
        _mystream_a15_source_stride_buf <= _mystream_a15_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_17 <= _mystream_a15_source_ram_rdata;
      end 
      if((_mystream_a15_source_fsm_15 == 1) && _mystream_stream_oready) begin
        _mystream_a15_idle <= 0;
        _mystream_a15_source_ram_raddr <= _mystream_a15_source_offset_buf;
        _mystream_a15_source_ram_renable <= 1;
        _mystream_a15_source_count <= _mystream_a15_source_size_buf;
      end 
      if((_mystream_a15_source_fsm_15 == 2) && _mystream_stream_oready) begin
        _mystream_a15_source_ram_raddr <= _mystream_a15_source_ram_raddr + _mystream_a15_source_stride_buf;
        _mystream_a15_source_ram_renable <= 1;
        _mystream_a15_source_count <= _mystream_a15_source_count - 1;
      end 
      if((_mystream_a15_source_fsm_15 == 2) && (_mystream_a15_source_count == 1) && _mystream_stream_oready) begin
        _mystream_a15_source_ram_renable <= 0;
        _mystream_a15_idle <= 1;
      end 
      if((_mystream_a15_source_fsm_15 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_a15_source_ram_renable <= 0;
        _mystream_a15_idle <= 1;
      end 
      if(_set_flag_233) begin
        _mystream_a16_source_mode <= 5'b1;
        _mystream_a16_source_offset <= _th_comp_offset_4;
        _mystream_a16_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_a16_source_stride <= 1;
      end 
      if(_set_flag_233) begin
        _mystream_a16_source_sel <= 17;
      end 
      if(_mystream_source_start && _mystream_a16_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_a16_source_offset_buf <= _mystream_a16_source_offset;
        _mystream_a16_source_size_buf <= _mystream_a16_source_size;
        _mystream_a16_source_stride_buf <= _mystream_a16_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_18 <= _mystream_a16_source_ram_rdata;
      end 
      if((_mystream_a16_source_fsm_16 == 1) && _mystream_stream_oready) begin
        _mystream_a16_idle <= 0;
        _mystream_a16_source_ram_raddr <= _mystream_a16_source_offset_buf;
        _mystream_a16_source_ram_renable <= 1;
        _mystream_a16_source_count <= _mystream_a16_source_size_buf;
      end 
      if((_mystream_a16_source_fsm_16 == 2) && _mystream_stream_oready) begin
        _mystream_a16_source_ram_raddr <= _mystream_a16_source_ram_raddr + _mystream_a16_source_stride_buf;
        _mystream_a16_source_ram_renable <= 1;
        _mystream_a16_source_count <= _mystream_a16_source_count - 1;
      end 
      if((_mystream_a16_source_fsm_16 == 2) && (_mystream_a16_source_count == 1) && _mystream_stream_oready) begin
        _mystream_a16_source_ram_renable <= 0;
        _mystream_a16_idle <= 1;
      end 
      if((_mystream_a16_source_fsm_16 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_a16_source_ram_renable <= 0;
        _mystream_a16_idle <= 1;
      end 
      if(_set_flag_236) begin
        _mystream_a17_source_mode <= 5'b1;
        _mystream_a17_source_offset <= _th_comp_offset_4;
        _mystream_a17_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_a17_source_stride <= 1;
      end 
      if(_set_flag_236) begin
        _mystream_a17_source_sel <= 18;
      end 
      if(_mystream_source_start && _mystream_a17_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_a17_source_offset_buf <= _mystream_a17_source_offset;
        _mystream_a17_source_size_buf <= _mystream_a17_source_size;
        _mystream_a17_source_stride_buf <= _mystream_a17_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_19 <= _mystream_a17_source_ram_rdata;
      end 
      if((_mystream_a17_source_fsm_17 == 1) && _mystream_stream_oready) begin
        _mystream_a17_idle <= 0;
        _mystream_a17_source_ram_raddr <= _mystream_a17_source_offset_buf;
        _mystream_a17_source_ram_renable <= 1;
        _mystream_a17_source_count <= _mystream_a17_source_size_buf;
      end 
      if((_mystream_a17_source_fsm_17 == 2) && _mystream_stream_oready) begin
        _mystream_a17_source_ram_raddr <= _mystream_a17_source_ram_raddr + _mystream_a17_source_stride_buf;
        _mystream_a17_source_ram_renable <= 1;
        _mystream_a17_source_count <= _mystream_a17_source_count - 1;
      end 
      if((_mystream_a17_source_fsm_17 == 2) && (_mystream_a17_source_count == 1) && _mystream_stream_oready) begin
        _mystream_a17_source_ram_renable <= 0;
        _mystream_a17_idle <= 1;
      end 
      if((_mystream_a17_source_fsm_17 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_a17_source_ram_renable <= 0;
        _mystream_a17_idle <= 1;
      end 
      if(_set_flag_239) begin
        _mystream_a18_source_mode <= 5'b1;
        _mystream_a18_source_offset <= _th_comp_offset_4;
        _mystream_a18_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_a18_source_stride <= 1;
      end 
      if(_set_flag_239) begin
        _mystream_a18_source_sel <= 19;
      end 
      if(_mystream_source_start && _mystream_a18_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_a18_source_offset_buf <= _mystream_a18_source_offset;
        _mystream_a18_source_size_buf <= _mystream_a18_source_size;
        _mystream_a18_source_stride_buf <= _mystream_a18_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_20 <= _mystream_a18_source_ram_rdata;
      end 
      if((_mystream_a18_source_fsm_18 == 1) && _mystream_stream_oready) begin
        _mystream_a18_idle <= 0;
        _mystream_a18_source_ram_raddr <= _mystream_a18_source_offset_buf;
        _mystream_a18_source_ram_renable <= 1;
        _mystream_a18_source_count <= _mystream_a18_source_size_buf;
      end 
      if((_mystream_a18_source_fsm_18 == 2) && _mystream_stream_oready) begin
        _mystream_a18_source_ram_raddr <= _mystream_a18_source_ram_raddr + _mystream_a18_source_stride_buf;
        _mystream_a18_source_ram_renable <= 1;
        _mystream_a18_source_count <= _mystream_a18_source_count - 1;
      end 
      if((_mystream_a18_source_fsm_18 == 2) && (_mystream_a18_source_count == 1) && _mystream_stream_oready) begin
        _mystream_a18_source_ram_renable <= 0;
        _mystream_a18_idle <= 1;
      end 
      if((_mystream_a18_source_fsm_18 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_a18_source_ram_renable <= 0;
        _mystream_a18_idle <= 1;
      end 
      if(_set_flag_242) begin
        _mystream_a19_source_mode <= 5'b1;
        _mystream_a19_source_offset <= _th_comp_offset_4;
        _mystream_a19_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_a19_source_stride <= 1;
      end 
      if(_set_flag_242) begin
        _mystream_a19_source_sel <= 20;
      end 
      if(_mystream_source_start && _mystream_a19_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_a19_source_offset_buf <= _mystream_a19_source_offset;
        _mystream_a19_source_size_buf <= _mystream_a19_source_size;
        _mystream_a19_source_stride_buf <= _mystream_a19_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_21 <= _mystream_a19_source_ram_rdata;
      end 
      if((_mystream_a19_source_fsm_19 == 1) && _mystream_stream_oready) begin
        _mystream_a19_idle <= 0;
        _mystream_a19_source_ram_raddr <= _mystream_a19_source_offset_buf;
        _mystream_a19_source_ram_renable <= 1;
        _mystream_a19_source_count <= _mystream_a19_source_size_buf;
      end 
      if((_mystream_a19_source_fsm_19 == 2) && _mystream_stream_oready) begin
        _mystream_a19_source_ram_raddr <= _mystream_a19_source_ram_raddr + _mystream_a19_source_stride_buf;
        _mystream_a19_source_ram_renable <= 1;
        _mystream_a19_source_count <= _mystream_a19_source_count - 1;
      end 
      if((_mystream_a19_source_fsm_19 == 2) && (_mystream_a19_source_count == 1) && _mystream_stream_oready) begin
        _mystream_a19_source_ram_renable <= 0;
        _mystream_a19_idle <= 1;
      end 
      if((_mystream_a19_source_fsm_19 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_a19_source_ram_renable <= 0;
        _mystream_a19_idle <= 1;
      end 
      if(_set_flag_245) begin
        _mystream_a20_source_mode <= 5'b1;
        _mystream_a20_source_offset <= _th_comp_offset_4;
        _mystream_a20_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_a20_source_stride <= 1;
      end 
      if(_set_flag_245) begin
        _mystream_a20_source_sel <= 21;
      end 
      if(_mystream_source_start && _mystream_a20_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_a20_source_offset_buf <= _mystream_a20_source_offset;
        _mystream_a20_source_size_buf <= _mystream_a20_source_size;
        _mystream_a20_source_stride_buf <= _mystream_a20_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_22 <= _mystream_a20_source_ram_rdata;
      end 
      if((_mystream_a20_source_fsm_20 == 1) && _mystream_stream_oready) begin
        _mystream_a20_idle <= 0;
        _mystream_a20_source_ram_raddr <= _mystream_a20_source_offset_buf;
        _mystream_a20_source_ram_renable <= 1;
        _mystream_a20_source_count <= _mystream_a20_source_size_buf;
      end 
      if((_mystream_a20_source_fsm_20 == 2) && _mystream_stream_oready) begin
        _mystream_a20_source_ram_raddr <= _mystream_a20_source_ram_raddr + _mystream_a20_source_stride_buf;
        _mystream_a20_source_ram_renable <= 1;
        _mystream_a20_source_count <= _mystream_a20_source_count - 1;
      end 
      if((_mystream_a20_source_fsm_20 == 2) && (_mystream_a20_source_count == 1) && _mystream_stream_oready) begin
        _mystream_a20_source_ram_renable <= 0;
        _mystream_a20_idle <= 1;
      end 
      if((_mystream_a20_source_fsm_20 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_a20_source_ram_renable <= 0;
        _mystream_a20_idle <= 1;
      end 
      if(_set_flag_248) begin
        _mystream_a21_source_mode <= 5'b1;
        _mystream_a21_source_offset <= _th_comp_offset_4;
        _mystream_a21_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_a21_source_stride <= 1;
      end 
      if(_set_flag_248) begin
        _mystream_a21_source_sel <= 22;
      end 
      if(_mystream_source_start && _mystream_a21_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_a21_source_offset_buf <= _mystream_a21_source_offset;
        _mystream_a21_source_size_buf <= _mystream_a21_source_size;
        _mystream_a21_source_stride_buf <= _mystream_a21_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_23 <= _mystream_a21_source_ram_rdata;
      end 
      if((_mystream_a21_source_fsm_21 == 1) && _mystream_stream_oready) begin
        _mystream_a21_idle <= 0;
        _mystream_a21_source_ram_raddr <= _mystream_a21_source_offset_buf;
        _mystream_a21_source_ram_renable <= 1;
        _mystream_a21_source_count <= _mystream_a21_source_size_buf;
      end 
      if((_mystream_a21_source_fsm_21 == 2) && _mystream_stream_oready) begin
        _mystream_a21_source_ram_raddr <= _mystream_a21_source_ram_raddr + _mystream_a21_source_stride_buf;
        _mystream_a21_source_ram_renable <= 1;
        _mystream_a21_source_count <= _mystream_a21_source_count - 1;
      end 
      if((_mystream_a21_source_fsm_21 == 2) && (_mystream_a21_source_count == 1) && _mystream_stream_oready) begin
        _mystream_a21_source_ram_renable <= 0;
        _mystream_a21_idle <= 1;
      end 
      if((_mystream_a21_source_fsm_21 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_a21_source_ram_renable <= 0;
        _mystream_a21_idle <= 1;
      end 
      if(_set_flag_251) begin
        _mystream_a22_source_mode <= 5'b1;
        _mystream_a22_source_offset <= _th_comp_offset_4;
        _mystream_a22_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_a22_source_stride <= 1;
      end 
      if(_set_flag_251) begin
        _mystream_a22_source_sel <= 23;
      end 
      if(_mystream_source_start && _mystream_a22_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_a22_source_offset_buf <= _mystream_a22_source_offset;
        _mystream_a22_source_size_buf <= _mystream_a22_source_size;
        _mystream_a22_source_stride_buf <= _mystream_a22_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_24 <= _mystream_a22_source_ram_rdata;
      end 
      if((_mystream_a22_source_fsm_22 == 1) && _mystream_stream_oready) begin
        _mystream_a22_idle <= 0;
        _mystream_a22_source_ram_raddr <= _mystream_a22_source_offset_buf;
        _mystream_a22_source_ram_renable <= 1;
        _mystream_a22_source_count <= _mystream_a22_source_size_buf;
      end 
      if((_mystream_a22_source_fsm_22 == 2) && _mystream_stream_oready) begin
        _mystream_a22_source_ram_raddr <= _mystream_a22_source_ram_raddr + _mystream_a22_source_stride_buf;
        _mystream_a22_source_ram_renable <= 1;
        _mystream_a22_source_count <= _mystream_a22_source_count - 1;
      end 
      if((_mystream_a22_source_fsm_22 == 2) && (_mystream_a22_source_count == 1) && _mystream_stream_oready) begin
        _mystream_a22_source_ram_renable <= 0;
        _mystream_a22_idle <= 1;
      end 
      if((_mystream_a22_source_fsm_22 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_a22_source_ram_renable <= 0;
        _mystream_a22_idle <= 1;
      end 
      if(_set_flag_254) begin
        _mystream_a23_source_mode <= 5'b1;
        _mystream_a23_source_offset <= _th_comp_offset_4;
        _mystream_a23_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_a23_source_stride <= 1;
      end 
      if(_set_flag_254) begin
        _mystream_a23_source_sel <= 24;
      end 
      if(_mystream_source_start && _mystream_a23_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_a23_source_offset_buf <= _mystream_a23_source_offset;
        _mystream_a23_source_size_buf <= _mystream_a23_source_size;
        _mystream_a23_source_stride_buf <= _mystream_a23_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_25 <= _mystream_a23_source_ram_rdata;
      end 
      if((_mystream_a23_source_fsm_23 == 1) && _mystream_stream_oready) begin
        _mystream_a23_idle <= 0;
        _mystream_a23_source_ram_raddr <= _mystream_a23_source_offset_buf;
        _mystream_a23_source_ram_renable <= 1;
        _mystream_a23_source_count <= _mystream_a23_source_size_buf;
      end 
      if((_mystream_a23_source_fsm_23 == 2) && _mystream_stream_oready) begin
        _mystream_a23_source_ram_raddr <= _mystream_a23_source_ram_raddr + _mystream_a23_source_stride_buf;
        _mystream_a23_source_ram_renable <= 1;
        _mystream_a23_source_count <= _mystream_a23_source_count - 1;
      end 
      if((_mystream_a23_source_fsm_23 == 2) && (_mystream_a23_source_count == 1) && _mystream_stream_oready) begin
        _mystream_a23_source_ram_renable <= 0;
        _mystream_a23_idle <= 1;
      end 
      if((_mystream_a23_source_fsm_23 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_a23_source_ram_renable <= 0;
        _mystream_a23_idle <= 1;
      end 
      if(_set_flag_257) begin
        _mystream_a24_source_mode <= 5'b1;
        _mystream_a24_source_offset <= _th_comp_offset_4;
        _mystream_a24_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_a24_source_stride <= 1;
      end 
      if(_set_flag_257) begin
        _mystream_a24_source_sel <= 25;
      end 
      if(_mystream_source_start && _mystream_a24_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_a24_source_offset_buf <= _mystream_a24_source_offset;
        _mystream_a24_source_size_buf <= _mystream_a24_source_size;
        _mystream_a24_source_stride_buf <= _mystream_a24_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_26 <= _mystream_a24_source_ram_rdata;
      end 
      if((_mystream_a24_source_fsm_24 == 1) && _mystream_stream_oready) begin
        _mystream_a24_idle <= 0;
        _mystream_a24_source_ram_raddr <= _mystream_a24_source_offset_buf;
        _mystream_a24_source_ram_renable <= 1;
        _mystream_a24_source_count <= _mystream_a24_source_size_buf;
      end 
      if((_mystream_a24_source_fsm_24 == 2) && _mystream_stream_oready) begin
        _mystream_a24_source_ram_raddr <= _mystream_a24_source_ram_raddr + _mystream_a24_source_stride_buf;
        _mystream_a24_source_ram_renable <= 1;
        _mystream_a24_source_count <= _mystream_a24_source_count - 1;
      end 
      if((_mystream_a24_source_fsm_24 == 2) && (_mystream_a24_source_count == 1) && _mystream_stream_oready) begin
        _mystream_a24_source_ram_renable <= 0;
        _mystream_a24_idle <= 1;
      end 
      if((_mystream_a24_source_fsm_24 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_a24_source_ram_renable <= 0;
        _mystream_a24_idle <= 1;
      end 
      if(_set_flag_260) begin
        _mystream_a25_source_mode <= 5'b1;
        _mystream_a25_source_offset <= _th_comp_offset_4;
        _mystream_a25_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_a25_source_stride <= 1;
      end 
      if(_set_flag_260) begin
        _mystream_a25_source_sel <= 26;
      end 
      if(_mystream_source_start && _mystream_a25_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_a25_source_offset_buf <= _mystream_a25_source_offset;
        _mystream_a25_source_size_buf <= _mystream_a25_source_size;
        _mystream_a25_source_stride_buf <= _mystream_a25_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_27 <= _mystream_a25_source_ram_rdata;
      end 
      if((_mystream_a25_source_fsm_25 == 1) && _mystream_stream_oready) begin
        _mystream_a25_idle <= 0;
        _mystream_a25_source_ram_raddr <= _mystream_a25_source_offset_buf;
        _mystream_a25_source_ram_renable <= 1;
        _mystream_a25_source_count <= _mystream_a25_source_size_buf;
      end 
      if((_mystream_a25_source_fsm_25 == 2) && _mystream_stream_oready) begin
        _mystream_a25_source_ram_raddr <= _mystream_a25_source_ram_raddr + _mystream_a25_source_stride_buf;
        _mystream_a25_source_ram_renable <= 1;
        _mystream_a25_source_count <= _mystream_a25_source_count - 1;
      end 
      if((_mystream_a25_source_fsm_25 == 2) && (_mystream_a25_source_count == 1) && _mystream_stream_oready) begin
        _mystream_a25_source_ram_renable <= 0;
        _mystream_a25_idle <= 1;
      end 
      if((_mystream_a25_source_fsm_25 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_a25_source_ram_renable <= 0;
        _mystream_a25_idle <= 1;
      end 
      if(_set_flag_263) begin
        _mystream_a26_source_mode <= 5'b1;
        _mystream_a26_source_offset <= _th_comp_offset_4;
        _mystream_a26_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_a26_source_stride <= 1;
      end 
      if(_set_flag_263) begin
        _mystream_a26_source_sel <= 27;
      end 
      if(_mystream_source_start && _mystream_a26_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_a26_source_offset_buf <= _mystream_a26_source_offset;
        _mystream_a26_source_size_buf <= _mystream_a26_source_size;
        _mystream_a26_source_stride_buf <= _mystream_a26_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_28 <= _mystream_a26_source_ram_rdata;
      end 
      if((_mystream_a26_source_fsm_26 == 1) && _mystream_stream_oready) begin
        _mystream_a26_idle <= 0;
        _mystream_a26_source_ram_raddr <= _mystream_a26_source_offset_buf;
        _mystream_a26_source_ram_renable <= 1;
        _mystream_a26_source_count <= _mystream_a26_source_size_buf;
      end 
      if((_mystream_a26_source_fsm_26 == 2) && _mystream_stream_oready) begin
        _mystream_a26_source_ram_raddr <= _mystream_a26_source_ram_raddr + _mystream_a26_source_stride_buf;
        _mystream_a26_source_ram_renable <= 1;
        _mystream_a26_source_count <= _mystream_a26_source_count - 1;
      end 
      if((_mystream_a26_source_fsm_26 == 2) && (_mystream_a26_source_count == 1) && _mystream_stream_oready) begin
        _mystream_a26_source_ram_renable <= 0;
        _mystream_a26_idle <= 1;
      end 
      if((_mystream_a26_source_fsm_26 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_a26_source_ram_renable <= 0;
        _mystream_a26_idle <= 1;
      end 
      if(_set_flag_266) begin
        _mystream_a27_source_mode <= 5'b1;
        _mystream_a27_source_offset <= _th_comp_offset_4;
        _mystream_a27_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_a27_source_stride <= 1;
      end 
      if(_set_flag_266) begin
        _mystream_a27_source_sel <= 28;
      end 
      if(_mystream_source_start && _mystream_a27_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_a27_source_offset_buf <= _mystream_a27_source_offset;
        _mystream_a27_source_size_buf <= _mystream_a27_source_size;
        _mystream_a27_source_stride_buf <= _mystream_a27_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_29 <= _mystream_a27_source_ram_rdata;
      end 
      if((_mystream_a27_source_fsm_27 == 1) && _mystream_stream_oready) begin
        _mystream_a27_idle <= 0;
        _mystream_a27_source_ram_raddr <= _mystream_a27_source_offset_buf;
        _mystream_a27_source_ram_renable <= 1;
        _mystream_a27_source_count <= _mystream_a27_source_size_buf;
      end 
      if((_mystream_a27_source_fsm_27 == 2) && _mystream_stream_oready) begin
        _mystream_a27_source_ram_raddr <= _mystream_a27_source_ram_raddr + _mystream_a27_source_stride_buf;
        _mystream_a27_source_ram_renable <= 1;
        _mystream_a27_source_count <= _mystream_a27_source_count - 1;
      end 
      if((_mystream_a27_source_fsm_27 == 2) && (_mystream_a27_source_count == 1) && _mystream_stream_oready) begin
        _mystream_a27_source_ram_renable <= 0;
        _mystream_a27_idle <= 1;
      end 
      if((_mystream_a27_source_fsm_27 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_a27_source_ram_renable <= 0;
        _mystream_a27_idle <= 1;
      end 
      if(_set_flag_269) begin
        _mystream_a28_source_mode <= 5'b1;
        _mystream_a28_source_offset <= _th_comp_offset_4;
        _mystream_a28_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_a28_source_stride <= 1;
      end 
      if(_set_flag_269) begin
        _mystream_a28_source_sel <= 29;
      end 
      if(_mystream_source_start && _mystream_a28_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_a28_source_offset_buf <= _mystream_a28_source_offset;
        _mystream_a28_source_size_buf <= _mystream_a28_source_size;
        _mystream_a28_source_stride_buf <= _mystream_a28_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_30 <= _mystream_a28_source_ram_rdata;
      end 
      if((_mystream_a28_source_fsm_28 == 1) && _mystream_stream_oready) begin
        _mystream_a28_idle <= 0;
        _mystream_a28_source_ram_raddr <= _mystream_a28_source_offset_buf;
        _mystream_a28_source_ram_renable <= 1;
        _mystream_a28_source_count <= _mystream_a28_source_size_buf;
      end 
      if((_mystream_a28_source_fsm_28 == 2) && _mystream_stream_oready) begin
        _mystream_a28_source_ram_raddr <= _mystream_a28_source_ram_raddr + _mystream_a28_source_stride_buf;
        _mystream_a28_source_ram_renable <= 1;
        _mystream_a28_source_count <= _mystream_a28_source_count - 1;
      end 
      if((_mystream_a28_source_fsm_28 == 2) && (_mystream_a28_source_count == 1) && _mystream_stream_oready) begin
        _mystream_a28_source_ram_renable <= 0;
        _mystream_a28_idle <= 1;
      end 
      if((_mystream_a28_source_fsm_28 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_a28_source_ram_renable <= 0;
        _mystream_a28_idle <= 1;
      end 
      if(_set_flag_272) begin
        _mystream_a29_source_mode <= 5'b1;
        _mystream_a29_source_offset <= _th_comp_offset_4;
        _mystream_a29_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_a29_source_stride <= 1;
      end 
      if(_set_flag_272) begin
        _mystream_a29_source_sel <= 30;
      end 
      if(_mystream_source_start && _mystream_a29_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_a29_source_offset_buf <= _mystream_a29_source_offset;
        _mystream_a29_source_size_buf <= _mystream_a29_source_size;
        _mystream_a29_source_stride_buf <= _mystream_a29_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_31 <= _mystream_a29_source_ram_rdata;
      end 
      if((_mystream_a29_source_fsm_29 == 1) && _mystream_stream_oready) begin
        _mystream_a29_idle <= 0;
        _mystream_a29_source_ram_raddr <= _mystream_a29_source_offset_buf;
        _mystream_a29_source_ram_renable <= 1;
        _mystream_a29_source_count <= _mystream_a29_source_size_buf;
      end 
      if((_mystream_a29_source_fsm_29 == 2) && _mystream_stream_oready) begin
        _mystream_a29_source_ram_raddr <= _mystream_a29_source_ram_raddr + _mystream_a29_source_stride_buf;
        _mystream_a29_source_ram_renable <= 1;
        _mystream_a29_source_count <= _mystream_a29_source_count - 1;
      end 
      if((_mystream_a29_source_fsm_29 == 2) && (_mystream_a29_source_count == 1) && _mystream_stream_oready) begin
        _mystream_a29_source_ram_renable <= 0;
        _mystream_a29_idle <= 1;
      end 
      if((_mystream_a29_source_fsm_29 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_a29_source_ram_renable <= 0;
        _mystream_a29_idle <= 1;
      end 
      if(_set_flag_275) begin
        _mystream_a30_source_mode <= 5'b1;
        _mystream_a30_source_offset <= _th_comp_offset_4;
        _mystream_a30_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_a30_source_stride <= 1;
      end 
      if(_set_flag_275) begin
        _mystream_a30_source_sel <= 31;
      end 
      if(_mystream_source_start && _mystream_a30_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_a30_source_offset_buf <= _mystream_a30_source_offset;
        _mystream_a30_source_size_buf <= _mystream_a30_source_size;
        _mystream_a30_source_stride_buf <= _mystream_a30_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_32 <= _mystream_a30_source_ram_rdata;
      end 
      if((_mystream_a30_source_fsm_30 == 1) && _mystream_stream_oready) begin
        _mystream_a30_idle <= 0;
        _mystream_a30_source_ram_raddr <= _mystream_a30_source_offset_buf;
        _mystream_a30_source_ram_renable <= 1;
        _mystream_a30_source_count <= _mystream_a30_source_size_buf;
      end 
      if((_mystream_a30_source_fsm_30 == 2) && _mystream_stream_oready) begin
        _mystream_a30_source_ram_raddr <= _mystream_a30_source_ram_raddr + _mystream_a30_source_stride_buf;
        _mystream_a30_source_ram_renable <= 1;
        _mystream_a30_source_count <= _mystream_a30_source_count - 1;
      end 
      if((_mystream_a30_source_fsm_30 == 2) && (_mystream_a30_source_count == 1) && _mystream_stream_oready) begin
        _mystream_a30_source_ram_renable <= 0;
        _mystream_a30_idle <= 1;
      end 
      if((_mystream_a30_source_fsm_30 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_a30_source_ram_renable <= 0;
        _mystream_a30_idle <= 1;
      end 
      if(_set_flag_278) begin
        _mystream_a31_source_mode <= 5'b1;
        _mystream_a31_source_offset <= _th_comp_offset_4;
        _mystream_a31_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_a31_source_stride <= 1;
      end 
      if(_set_flag_278) begin
        _mystream_a31_source_sel <= 32;
      end 
      if(_mystream_source_start && _mystream_a31_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_a31_source_offset_buf <= _mystream_a31_source_offset;
        _mystream_a31_source_size_buf <= _mystream_a31_source_size;
        _mystream_a31_source_stride_buf <= _mystream_a31_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_33 <= _mystream_a31_source_ram_rdata;
      end 
      if((_mystream_a31_source_fsm_31 == 1) && _mystream_stream_oready) begin
        _mystream_a31_idle <= 0;
        _mystream_a31_source_ram_raddr <= _mystream_a31_source_offset_buf;
        _mystream_a31_source_ram_renable <= 1;
        _mystream_a31_source_count <= _mystream_a31_source_size_buf;
      end 
      if((_mystream_a31_source_fsm_31 == 2) && _mystream_stream_oready) begin
        _mystream_a31_source_ram_raddr <= _mystream_a31_source_ram_raddr + _mystream_a31_source_stride_buf;
        _mystream_a31_source_ram_renable <= 1;
        _mystream_a31_source_count <= _mystream_a31_source_count - 1;
      end 
      if((_mystream_a31_source_fsm_31 == 2) && (_mystream_a31_source_count == 1) && _mystream_stream_oready) begin
        _mystream_a31_source_ram_renable <= 0;
        _mystream_a31_idle <= 1;
      end 
      if((_mystream_a31_source_fsm_31 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_a31_source_ram_renable <= 0;
        _mystream_a31_idle <= 1;
      end 
      if(_set_flag_281) begin
        _mystream_b0_source_mode <= 5'b1;
        _mystream_b0_source_offset <= _th_comp_offset_4;
        _mystream_b0_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_b0_source_stride <= 1;
      end 
      if(_set_flag_281) begin
        _mystream_b0_source_sel <= 33;
      end 
      if(_mystream_source_start && _mystream_b0_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_b0_source_offset_buf <= _mystream_b0_source_offset;
        _mystream_b0_source_size_buf <= _mystream_b0_source_size;
        _mystream_b0_source_stride_buf <= _mystream_b0_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_34 <= _mystream_b0_source_ram_rdata;
      end 
      if((_mystream_b0_source_fsm_32 == 1) && _mystream_stream_oready) begin
        _mystream_b0_idle <= 0;
        _mystream_b0_source_ram_raddr <= _mystream_b0_source_offset_buf;
        _mystream_b0_source_ram_renable <= 1;
        _mystream_b0_source_count <= _mystream_b0_source_size_buf;
      end 
      if((_mystream_b0_source_fsm_32 == 2) && _mystream_stream_oready) begin
        _mystream_b0_source_ram_raddr <= _mystream_b0_source_ram_raddr + _mystream_b0_source_stride_buf;
        _mystream_b0_source_ram_renable <= 1;
        _mystream_b0_source_count <= _mystream_b0_source_count - 1;
      end 
      if((_mystream_b0_source_fsm_32 == 2) && (_mystream_b0_source_count == 1) && _mystream_stream_oready) begin
        _mystream_b0_source_ram_renable <= 0;
        _mystream_b0_idle <= 1;
      end 
      if((_mystream_b0_source_fsm_32 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_b0_source_ram_renable <= 0;
        _mystream_b0_idle <= 1;
      end 
      if(_set_flag_284) begin
        _mystream_b1_source_mode <= 5'b1;
        _mystream_b1_source_offset <= _th_comp_offset_4;
        _mystream_b1_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_b1_source_stride <= 1;
      end 
      if(_set_flag_284) begin
        _mystream_b1_source_sel <= 34;
      end 
      if(_mystream_source_start && _mystream_b1_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_b1_source_offset_buf <= _mystream_b1_source_offset;
        _mystream_b1_source_size_buf <= _mystream_b1_source_size;
        _mystream_b1_source_stride_buf <= _mystream_b1_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_35 <= _mystream_b1_source_ram_rdata;
      end 
      if((_mystream_b1_source_fsm_33 == 1) && _mystream_stream_oready) begin
        _mystream_b1_idle <= 0;
        _mystream_b1_source_ram_raddr <= _mystream_b1_source_offset_buf;
        _mystream_b1_source_ram_renable <= 1;
        _mystream_b1_source_count <= _mystream_b1_source_size_buf;
      end 
      if((_mystream_b1_source_fsm_33 == 2) && _mystream_stream_oready) begin
        _mystream_b1_source_ram_raddr <= _mystream_b1_source_ram_raddr + _mystream_b1_source_stride_buf;
        _mystream_b1_source_ram_renable <= 1;
        _mystream_b1_source_count <= _mystream_b1_source_count - 1;
      end 
      if((_mystream_b1_source_fsm_33 == 2) && (_mystream_b1_source_count == 1) && _mystream_stream_oready) begin
        _mystream_b1_source_ram_renable <= 0;
        _mystream_b1_idle <= 1;
      end 
      if((_mystream_b1_source_fsm_33 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_b1_source_ram_renable <= 0;
        _mystream_b1_idle <= 1;
      end 
      if(_set_flag_287) begin
        _mystream_b2_source_mode <= 5'b1;
        _mystream_b2_source_offset <= _th_comp_offset_4;
        _mystream_b2_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_b2_source_stride <= 1;
      end 
      if(_set_flag_287) begin
        _mystream_b2_source_sel <= 35;
      end 
      if(_mystream_source_start && _mystream_b2_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_b2_source_offset_buf <= _mystream_b2_source_offset;
        _mystream_b2_source_size_buf <= _mystream_b2_source_size;
        _mystream_b2_source_stride_buf <= _mystream_b2_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_36 <= _mystream_b2_source_ram_rdata;
      end 
      if((_mystream_b2_source_fsm_34 == 1) && _mystream_stream_oready) begin
        _mystream_b2_idle <= 0;
        _mystream_b2_source_ram_raddr <= _mystream_b2_source_offset_buf;
        _mystream_b2_source_ram_renable <= 1;
        _mystream_b2_source_count <= _mystream_b2_source_size_buf;
      end 
      if((_mystream_b2_source_fsm_34 == 2) && _mystream_stream_oready) begin
        _mystream_b2_source_ram_raddr <= _mystream_b2_source_ram_raddr + _mystream_b2_source_stride_buf;
        _mystream_b2_source_ram_renable <= 1;
        _mystream_b2_source_count <= _mystream_b2_source_count - 1;
      end 
      if((_mystream_b2_source_fsm_34 == 2) && (_mystream_b2_source_count == 1) && _mystream_stream_oready) begin
        _mystream_b2_source_ram_renable <= 0;
        _mystream_b2_idle <= 1;
      end 
      if((_mystream_b2_source_fsm_34 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_b2_source_ram_renable <= 0;
        _mystream_b2_idle <= 1;
      end 
      if(_set_flag_290) begin
        _mystream_b3_source_mode <= 5'b1;
        _mystream_b3_source_offset <= _th_comp_offset_4;
        _mystream_b3_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_b3_source_stride <= 1;
      end 
      if(_set_flag_290) begin
        _mystream_b3_source_sel <= 36;
      end 
      if(_mystream_source_start && _mystream_b3_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_b3_source_offset_buf <= _mystream_b3_source_offset;
        _mystream_b3_source_size_buf <= _mystream_b3_source_size;
        _mystream_b3_source_stride_buf <= _mystream_b3_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_37 <= _mystream_b3_source_ram_rdata;
      end 
      if((_mystream_b3_source_fsm_35 == 1) && _mystream_stream_oready) begin
        _mystream_b3_idle <= 0;
        _mystream_b3_source_ram_raddr <= _mystream_b3_source_offset_buf;
        _mystream_b3_source_ram_renable <= 1;
        _mystream_b3_source_count <= _mystream_b3_source_size_buf;
      end 
      if((_mystream_b3_source_fsm_35 == 2) && _mystream_stream_oready) begin
        _mystream_b3_source_ram_raddr <= _mystream_b3_source_ram_raddr + _mystream_b3_source_stride_buf;
        _mystream_b3_source_ram_renable <= 1;
        _mystream_b3_source_count <= _mystream_b3_source_count - 1;
      end 
      if((_mystream_b3_source_fsm_35 == 2) && (_mystream_b3_source_count == 1) && _mystream_stream_oready) begin
        _mystream_b3_source_ram_renable <= 0;
        _mystream_b3_idle <= 1;
      end 
      if((_mystream_b3_source_fsm_35 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_b3_source_ram_renable <= 0;
        _mystream_b3_idle <= 1;
      end 
      if(_set_flag_293) begin
        _mystream_b4_source_mode <= 5'b1;
        _mystream_b4_source_offset <= _th_comp_offset_4;
        _mystream_b4_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_b4_source_stride <= 1;
      end 
      if(_set_flag_293) begin
        _mystream_b4_source_sel <= 37;
      end 
      if(_mystream_source_start && _mystream_b4_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_b4_source_offset_buf <= _mystream_b4_source_offset;
        _mystream_b4_source_size_buf <= _mystream_b4_source_size;
        _mystream_b4_source_stride_buf <= _mystream_b4_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_38 <= _mystream_b4_source_ram_rdata;
      end 
      if((_mystream_b4_source_fsm_36 == 1) && _mystream_stream_oready) begin
        _mystream_b4_idle <= 0;
        _mystream_b4_source_ram_raddr <= _mystream_b4_source_offset_buf;
        _mystream_b4_source_ram_renable <= 1;
        _mystream_b4_source_count <= _mystream_b4_source_size_buf;
      end 
      if((_mystream_b4_source_fsm_36 == 2) && _mystream_stream_oready) begin
        _mystream_b4_source_ram_raddr <= _mystream_b4_source_ram_raddr + _mystream_b4_source_stride_buf;
        _mystream_b4_source_ram_renable <= 1;
        _mystream_b4_source_count <= _mystream_b4_source_count - 1;
      end 
      if((_mystream_b4_source_fsm_36 == 2) && (_mystream_b4_source_count == 1) && _mystream_stream_oready) begin
        _mystream_b4_source_ram_renable <= 0;
        _mystream_b4_idle <= 1;
      end 
      if((_mystream_b4_source_fsm_36 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_b4_source_ram_renable <= 0;
        _mystream_b4_idle <= 1;
      end 
      if(_set_flag_296) begin
        _mystream_b5_source_mode <= 5'b1;
        _mystream_b5_source_offset <= _th_comp_offset_4;
        _mystream_b5_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_b5_source_stride <= 1;
      end 
      if(_set_flag_296) begin
        _mystream_b5_source_sel <= 38;
      end 
      if(_mystream_source_start && _mystream_b5_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_b5_source_offset_buf <= _mystream_b5_source_offset;
        _mystream_b5_source_size_buf <= _mystream_b5_source_size;
        _mystream_b5_source_stride_buf <= _mystream_b5_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_39 <= _mystream_b5_source_ram_rdata;
      end 
      if((_mystream_b5_source_fsm_37 == 1) && _mystream_stream_oready) begin
        _mystream_b5_idle <= 0;
        _mystream_b5_source_ram_raddr <= _mystream_b5_source_offset_buf;
        _mystream_b5_source_ram_renable <= 1;
        _mystream_b5_source_count <= _mystream_b5_source_size_buf;
      end 
      if((_mystream_b5_source_fsm_37 == 2) && _mystream_stream_oready) begin
        _mystream_b5_source_ram_raddr <= _mystream_b5_source_ram_raddr + _mystream_b5_source_stride_buf;
        _mystream_b5_source_ram_renable <= 1;
        _mystream_b5_source_count <= _mystream_b5_source_count - 1;
      end 
      if((_mystream_b5_source_fsm_37 == 2) && (_mystream_b5_source_count == 1) && _mystream_stream_oready) begin
        _mystream_b5_source_ram_renable <= 0;
        _mystream_b5_idle <= 1;
      end 
      if((_mystream_b5_source_fsm_37 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_b5_source_ram_renable <= 0;
        _mystream_b5_idle <= 1;
      end 
      if(_set_flag_299) begin
        _mystream_b6_source_mode <= 5'b1;
        _mystream_b6_source_offset <= _th_comp_offset_4;
        _mystream_b6_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_b6_source_stride <= 1;
      end 
      if(_set_flag_299) begin
        _mystream_b6_source_sel <= 39;
      end 
      if(_mystream_source_start && _mystream_b6_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_b6_source_offset_buf <= _mystream_b6_source_offset;
        _mystream_b6_source_size_buf <= _mystream_b6_source_size;
        _mystream_b6_source_stride_buf <= _mystream_b6_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_40 <= _mystream_b6_source_ram_rdata;
      end 
      if((_mystream_b6_source_fsm_38 == 1) && _mystream_stream_oready) begin
        _mystream_b6_idle <= 0;
        _mystream_b6_source_ram_raddr <= _mystream_b6_source_offset_buf;
        _mystream_b6_source_ram_renable <= 1;
        _mystream_b6_source_count <= _mystream_b6_source_size_buf;
      end 
      if((_mystream_b6_source_fsm_38 == 2) && _mystream_stream_oready) begin
        _mystream_b6_source_ram_raddr <= _mystream_b6_source_ram_raddr + _mystream_b6_source_stride_buf;
        _mystream_b6_source_ram_renable <= 1;
        _mystream_b6_source_count <= _mystream_b6_source_count - 1;
      end 
      if((_mystream_b6_source_fsm_38 == 2) && (_mystream_b6_source_count == 1) && _mystream_stream_oready) begin
        _mystream_b6_source_ram_renable <= 0;
        _mystream_b6_idle <= 1;
      end 
      if((_mystream_b6_source_fsm_38 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_b6_source_ram_renable <= 0;
        _mystream_b6_idle <= 1;
      end 
      if(_set_flag_302) begin
        _mystream_b7_source_mode <= 5'b1;
        _mystream_b7_source_offset <= _th_comp_offset_4;
        _mystream_b7_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_b7_source_stride <= 1;
      end 
      if(_set_flag_302) begin
        _mystream_b7_source_sel <= 40;
      end 
      if(_mystream_source_start && _mystream_b7_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_b7_source_offset_buf <= _mystream_b7_source_offset;
        _mystream_b7_source_size_buf <= _mystream_b7_source_size;
        _mystream_b7_source_stride_buf <= _mystream_b7_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_41 <= _mystream_b7_source_ram_rdata;
      end 
      if((_mystream_b7_source_fsm_39 == 1) && _mystream_stream_oready) begin
        _mystream_b7_idle <= 0;
        _mystream_b7_source_ram_raddr <= _mystream_b7_source_offset_buf;
        _mystream_b7_source_ram_renable <= 1;
        _mystream_b7_source_count <= _mystream_b7_source_size_buf;
      end 
      if((_mystream_b7_source_fsm_39 == 2) && _mystream_stream_oready) begin
        _mystream_b7_source_ram_raddr <= _mystream_b7_source_ram_raddr + _mystream_b7_source_stride_buf;
        _mystream_b7_source_ram_renable <= 1;
        _mystream_b7_source_count <= _mystream_b7_source_count - 1;
      end 
      if((_mystream_b7_source_fsm_39 == 2) && (_mystream_b7_source_count == 1) && _mystream_stream_oready) begin
        _mystream_b7_source_ram_renable <= 0;
        _mystream_b7_idle <= 1;
      end 
      if((_mystream_b7_source_fsm_39 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_b7_source_ram_renable <= 0;
        _mystream_b7_idle <= 1;
      end 
      if(_set_flag_305) begin
        _mystream_b8_source_mode <= 5'b1;
        _mystream_b8_source_offset <= _th_comp_offset_4;
        _mystream_b8_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_b8_source_stride <= 1;
      end 
      if(_set_flag_305) begin
        _mystream_b8_source_sel <= 41;
      end 
      if(_mystream_source_start && _mystream_b8_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_b8_source_offset_buf <= _mystream_b8_source_offset;
        _mystream_b8_source_size_buf <= _mystream_b8_source_size;
        _mystream_b8_source_stride_buf <= _mystream_b8_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_42 <= _mystream_b8_source_ram_rdata;
      end 
      if((_mystream_b8_source_fsm_40 == 1) && _mystream_stream_oready) begin
        _mystream_b8_idle <= 0;
        _mystream_b8_source_ram_raddr <= _mystream_b8_source_offset_buf;
        _mystream_b8_source_ram_renable <= 1;
        _mystream_b8_source_count <= _mystream_b8_source_size_buf;
      end 
      if((_mystream_b8_source_fsm_40 == 2) && _mystream_stream_oready) begin
        _mystream_b8_source_ram_raddr <= _mystream_b8_source_ram_raddr + _mystream_b8_source_stride_buf;
        _mystream_b8_source_ram_renable <= 1;
        _mystream_b8_source_count <= _mystream_b8_source_count - 1;
      end 
      if((_mystream_b8_source_fsm_40 == 2) && (_mystream_b8_source_count == 1) && _mystream_stream_oready) begin
        _mystream_b8_source_ram_renable <= 0;
        _mystream_b8_idle <= 1;
      end 
      if((_mystream_b8_source_fsm_40 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_b8_source_ram_renable <= 0;
        _mystream_b8_idle <= 1;
      end 
      if(_set_flag_308) begin
        _mystream_b9_source_mode <= 5'b1;
        _mystream_b9_source_offset <= _th_comp_offset_4;
        _mystream_b9_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_b9_source_stride <= 1;
      end 
      if(_set_flag_308) begin
        _mystream_b9_source_sel <= 42;
      end 
      if(_mystream_source_start && _mystream_b9_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_b9_source_offset_buf <= _mystream_b9_source_offset;
        _mystream_b9_source_size_buf <= _mystream_b9_source_size;
        _mystream_b9_source_stride_buf <= _mystream_b9_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_43 <= _mystream_b9_source_ram_rdata;
      end 
      if((_mystream_b9_source_fsm_41 == 1) && _mystream_stream_oready) begin
        _mystream_b9_idle <= 0;
        _mystream_b9_source_ram_raddr <= _mystream_b9_source_offset_buf;
        _mystream_b9_source_ram_renable <= 1;
        _mystream_b9_source_count <= _mystream_b9_source_size_buf;
      end 
      if((_mystream_b9_source_fsm_41 == 2) && _mystream_stream_oready) begin
        _mystream_b9_source_ram_raddr <= _mystream_b9_source_ram_raddr + _mystream_b9_source_stride_buf;
        _mystream_b9_source_ram_renable <= 1;
        _mystream_b9_source_count <= _mystream_b9_source_count - 1;
      end 
      if((_mystream_b9_source_fsm_41 == 2) && (_mystream_b9_source_count == 1) && _mystream_stream_oready) begin
        _mystream_b9_source_ram_renable <= 0;
        _mystream_b9_idle <= 1;
      end 
      if((_mystream_b9_source_fsm_41 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_b9_source_ram_renable <= 0;
        _mystream_b9_idle <= 1;
      end 
      if(_set_flag_311) begin
        _mystream_b10_source_mode <= 5'b1;
        _mystream_b10_source_offset <= _th_comp_offset_4;
        _mystream_b10_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_b10_source_stride <= 1;
      end 
      if(_set_flag_311) begin
        _mystream_b10_source_sel <= 43;
      end 
      if(_mystream_source_start && _mystream_b10_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_b10_source_offset_buf <= _mystream_b10_source_offset;
        _mystream_b10_source_size_buf <= _mystream_b10_source_size;
        _mystream_b10_source_stride_buf <= _mystream_b10_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_44 <= _mystream_b10_source_ram_rdata;
      end 
      if((_mystream_b10_source_fsm_42 == 1) && _mystream_stream_oready) begin
        _mystream_b10_idle <= 0;
        _mystream_b10_source_ram_raddr <= _mystream_b10_source_offset_buf;
        _mystream_b10_source_ram_renable <= 1;
        _mystream_b10_source_count <= _mystream_b10_source_size_buf;
      end 
      if((_mystream_b10_source_fsm_42 == 2) && _mystream_stream_oready) begin
        _mystream_b10_source_ram_raddr <= _mystream_b10_source_ram_raddr + _mystream_b10_source_stride_buf;
        _mystream_b10_source_ram_renable <= 1;
        _mystream_b10_source_count <= _mystream_b10_source_count - 1;
      end 
      if((_mystream_b10_source_fsm_42 == 2) && (_mystream_b10_source_count == 1) && _mystream_stream_oready) begin
        _mystream_b10_source_ram_renable <= 0;
        _mystream_b10_idle <= 1;
      end 
      if((_mystream_b10_source_fsm_42 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_b10_source_ram_renable <= 0;
        _mystream_b10_idle <= 1;
      end 
      if(_set_flag_314) begin
        _mystream_b11_source_mode <= 5'b1;
        _mystream_b11_source_offset <= _th_comp_offset_4;
        _mystream_b11_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_b11_source_stride <= 1;
      end 
      if(_set_flag_314) begin
        _mystream_b11_source_sel <= 44;
      end 
      if(_mystream_source_start && _mystream_b11_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_b11_source_offset_buf <= _mystream_b11_source_offset;
        _mystream_b11_source_size_buf <= _mystream_b11_source_size;
        _mystream_b11_source_stride_buf <= _mystream_b11_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_45 <= _mystream_b11_source_ram_rdata;
      end 
      if((_mystream_b11_source_fsm_43 == 1) && _mystream_stream_oready) begin
        _mystream_b11_idle <= 0;
        _mystream_b11_source_ram_raddr <= _mystream_b11_source_offset_buf;
        _mystream_b11_source_ram_renable <= 1;
        _mystream_b11_source_count <= _mystream_b11_source_size_buf;
      end 
      if((_mystream_b11_source_fsm_43 == 2) && _mystream_stream_oready) begin
        _mystream_b11_source_ram_raddr <= _mystream_b11_source_ram_raddr + _mystream_b11_source_stride_buf;
        _mystream_b11_source_ram_renable <= 1;
        _mystream_b11_source_count <= _mystream_b11_source_count - 1;
      end 
      if((_mystream_b11_source_fsm_43 == 2) && (_mystream_b11_source_count == 1) && _mystream_stream_oready) begin
        _mystream_b11_source_ram_renable <= 0;
        _mystream_b11_idle <= 1;
      end 
      if((_mystream_b11_source_fsm_43 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_b11_source_ram_renable <= 0;
        _mystream_b11_idle <= 1;
      end 
      if(_set_flag_317) begin
        _mystream_b12_source_mode <= 5'b1;
        _mystream_b12_source_offset <= _th_comp_offset_4;
        _mystream_b12_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_b12_source_stride <= 1;
      end 
      if(_set_flag_317) begin
        _mystream_b12_source_sel <= 45;
      end 
      if(_mystream_source_start && _mystream_b12_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_b12_source_offset_buf <= _mystream_b12_source_offset;
        _mystream_b12_source_size_buf <= _mystream_b12_source_size;
        _mystream_b12_source_stride_buf <= _mystream_b12_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_46 <= _mystream_b12_source_ram_rdata;
      end 
      if((_mystream_b12_source_fsm_44 == 1) && _mystream_stream_oready) begin
        _mystream_b12_idle <= 0;
        _mystream_b12_source_ram_raddr <= _mystream_b12_source_offset_buf;
        _mystream_b12_source_ram_renable <= 1;
        _mystream_b12_source_count <= _mystream_b12_source_size_buf;
      end 
      if((_mystream_b12_source_fsm_44 == 2) && _mystream_stream_oready) begin
        _mystream_b12_source_ram_raddr <= _mystream_b12_source_ram_raddr + _mystream_b12_source_stride_buf;
        _mystream_b12_source_ram_renable <= 1;
        _mystream_b12_source_count <= _mystream_b12_source_count - 1;
      end 
      if((_mystream_b12_source_fsm_44 == 2) && (_mystream_b12_source_count == 1) && _mystream_stream_oready) begin
        _mystream_b12_source_ram_renable <= 0;
        _mystream_b12_idle <= 1;
      end 
      if((_mystream_b12_source_fsm_44 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_b12_source_ram_renable <= 0;
        _mystream_b12_idle <= 1;
      end 
      if(_set_flag_320) begin
        _mystream_b13_source_mode <= 5'b1;
        _mystream_b13_source_offset <= _th_comp_offset_4;
        _mystream_b13_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_b13_source_stride <= 1;
      end 
      if(_set_flag_320) begin
        _mystream_b13_source_sel <= 46;
      end 
      if(_mystream_source_start && _mystream_b13_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_b13_source_offset_buf <= _mystream_b13_source_offset;
        _mystream_b13_source_size_buf <= _mystream_b13_source_size;
        _mystream_b13_source_stride_buf <= _mystream_b13_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_47 <= _mystream_b13_source_ram_rdata;
      end 
      if((_mystream_b13_source_fsm_45 == 1) && _mystream_stream_oready) begin
        _mystream_b13_idle <= 0;
        _mystream_b13_source_ram_raddr <= _mystream_b13_source_offset_buf;
        _mystream_b13_source_ram_renable <= 1;
        _mystream_b13_source_count <= _mystream_b13_source_size_buf;
      end 
      if((_mystream_b13_source_fsm_45 == 2) && _mystream_stream_oready) begin
        _mystream_b13_source_ram_raddr <= _mystream_b13_source_ram_raddr + _mystream_b13_source_stride_buf;
        _mystream_b13_source_ram_renable <= 1;
        _mystream_b13_source_count <= _mystream_b13_source_count - 1;
      end 
      if((_mystream_b13_source_fsm_45 == 2) && (_mystream_b13_source_count == 1) && _mystream_stream_oready) begin
        _mystream_b13_source_ram_renable <= 0;
        _mystream_b13_idle <= 1;
      end 
      if((_mystream_b13_source_fsm_45 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_b13_source_ram_renable <= 0;
        _mystream_b13_idle <= 1;
      end 
      if(_set_flag_323) begin
        _mystream_b14_source_mode <= 5'b1;
        _mystream_b14_source_offset <= _th_comp_offset_4;
        _mystream_b14_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_b14_source_stride <= 1;
      end 
      if(_set_flag_323) begin
        _mystream_b14_source_sel <= 47;
      end 
      if(_mystream_source_start && _mystream_b14_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_b14_source_offset_buf <= _mystream_b14_source_offset;
        _mystream_b14_source_size_buf <= _mystream_b14_source_size;
        _mystream_b14_source_stride_buf <= _mystream_b14_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_48 <= _mystream_b14_source_ram_rdata;
      end 
      if((_mystream_b14_source_fsm_46 == 1) && _mystream_stream_oready) begin
        _mystream_b14_idle <= 0;
        _mystream_b14_source_ram_raddr <= _mystream_b14_source_offset_buf;
        _mystream_b14_source_ram_renable <= 1;
        _mystream_b14_source_count <= _mystream_b14_source_size_buf;
      end 
      if((_mystream_b14_source_fsm_46 == 2) && _mystream_stream_oready) begin
        _mystream_b14_source_ram_raddr <= _mystream_b14_source_ram_raddr + _mystream_b14_source_stride_buf;
        _mystream_b14_source_ram_renable <= 1;
        _mystream_b14_source_count <= _mystream_b14_source_count - 1;
      end 
      if((_mystream_b14_source_fsm_46 == 2) && (_mystream_b14_source_count == 1) && _mystream_stream_oready) begin
        _mystream_b14_source_ram_renable <= 0;
        _mystream_b14_idle <= 1;
      end 
      if((_mystream_b14_source_fsm_46 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_b14_source_ram_renable <= 0;
        _mystream_b14_idle <= 1;
      end 
      if(_set_flag_326) begin
        _mystream_b15_source_mode <= 5'b1;
        _mystream_b15_source_offset <= _th_comp_offset_4;
        _mystream_b15_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_b15_source_stride <= 1;
      end 
      if(_set_flag_326) begin
        _mystream_b15_source_sel <= 48;
      end 
      if(_mystream_source_start && _mystream_b15_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_b15_source_offset_buf <= _mystream_b15_source_offset;
        _mystream_b15_source_size_buf <= _mystream_b15_source_size;
        _mystream_b15_source_stride_buf <= _mystream_b15_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_49 <= _mystream_b15_source_ram_rdata;
      end 
      if((_mystream_b15_source_fsm_47 == 1) && _mystream_stream_oready) begin
        _mystream_b15_idle <= 0;
        _mystream_b15_source_ram_raddr <= _mystream_b15_source_offset_buf;
        _mystream_b15_source_ram_renable <= 1;
        _mystream_b15_source_count <= _mystream_b15_source_size_buf;
      end 
      if((_mystream_b15_source_fsm_47 == 2) && _mystream_stream_oready) begin
        _mystream_b15_source_ram_raddr <= _mystream_b15_source_ram_raddr + _mystream_b15_source_stride_buf;
        _mystream_b15_source_ram_renable <= 1;
        _mystream_b15_source_count <= _mystream_b15_source_count - 1;
      end 
      if((_mystream_b15_source_fsm_47 == 2) && (_mystream_b15_source_count == 1) && _mystream_stream_oready) begin
        _mystream_b15_source_ram_renable <= 0;
        _mystream_b15_idle <= 1;
      end 
      if((_mystream_b15_source_fsm_47 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_b15_source_ram_renable <= 0;
        _mystream_b15_idle <= 1;
      end 
      if(_set_flag_329) begin
        _mystream_b16_source_mode <= 5'b1;
        _mystream_b16_source_offset <= _th_comp_offset_4;
        _mystream_b16_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_b16_source_stride <= 1;
      end 
      if(_set_flag_329) begin
        _mystream_b16_source_sel <= 49;
      end 
      if(_mystream_source_start && _mystream_b16_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_b16_source_offset_buf <= _mystream_b16_source_offset;
        _mystream_b16_source_size_buf <= _mystream_b16_source_size;
        _mystream_b16_source_stride_buf <= _mystream_b16_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_50 <= _mystream_b16_source_ram_rdata;
      end 
      if((_mystream_b16_source_fsm_48 == 1) && _mystream_stream_oready) begin
        _mystream_b16_idle <= 0;
        _mystream_b16_source_ram_raddr <= _mystream_b16_source_offset_buf;
        _mystream_b16_source_ram_renable <= 1;
        _mystream_b16_source_count <= _mystream_b16_source_size_buf;
      end 
      if((_mystream_b16_source_fsm_48 == 2) && _mystream_stream_oready) begin
        _mystream_b16_source_ram_raddr <= _mystream_b16_source_ram_raddr + _mystream_b16_source_stride_buf;
        _mystream_b16_source_ram_renable <= 1;
        _mystream_b16_source_count <= _mystream_b16_source_count - 1;
      end 
      if((_mystream_b16_source_fsm_48 == 2) && (_mystream_b16_source_count == 1) && _mystream_stream_oready) begin
        _mystream_b16_source_ram_renable <= 0;
        _mystream_b16_idle <= 1;
      end 
      if((_mystream_b16_source_fsm_48 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_b16_source_ram_renable <= 0;
        _mystream_b16_idle <= 1;
      end 
      if(_set_flag_332) begin
        _mystream_b17_source_mode <= 5'b1;
        _mystream_b17_source_offset <= _th_comp_offset_4;
        _mystream_b17_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_b17_source_stride <= 1;
      end 
      if(_set_flag_332) begin
        _mystream_b17_source_sel <= 50;
      end 
      if(_mystream_source_start && _mystream_b17_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_b17_source_offset_buf <= _mystream_b17_source_offset;
        _mystream_b17_source_size_buf <= _mystream_b17_source_size;
        _mystream_b17_source_stride_buf <= _mystream_b17_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_51 <= _mystream_b17_source_ram_rdata;
      end 
      if((_mystream_b17_source_fsm_49 == 1) && _mystream_stream_oready) begin
        _mystream_b17_idle <= 0;
        _mystream_b17_source_ram_raddr <= _mystream_b17_source_offset_buf;
        _mystream_b17_source_ram_renable <= 1;
        _mystream_b17_source_count <= _mystream_b17_source_size_buf;
      end 
      if((_mystream_b17_source_fsm_49 == 2) && _mystream_stream_oready) begin
        _mystream_b17_source_ram_raddr <= _mystream_b17_source_ram_raddr + _mystream_b17_source_stride_buf;
        _mystream_b17_source_ram_renable <= 1;
        _mystream_b17_source_count <= _mystream_b17_source_count - 1;
      end 
      if((_mystream_b17_source_fsm_49 == 2) && (_mystream_b17_source_count == 1) && _mystream_stream_oready) begin
        _mystream_b17_source_ram_renable <= 0;
        _mystream_b17_idle <= 1;
      end 
      if((_mystream_b17_source_fsm_49 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_b17_source_ram_renable <= 0;
        _mystream_b17_idle <= 1;
      end 
      if(_set_flag_335) begin
        _mystream_b18_source_mode <= 5'b1;
        _mystream_b18_source_offset <= _th_comp_offset_4;
        _mystream_b18_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_b18_source_stride <= 1;
      end 
      if(_set_flag_335) begin
        _mystream_b18_source_sel <= 51;
      end 
      if(_mystream_source_start && _mystream_b18_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_b18_source_offset_buf <= _mystream_b18_source_offset;
        _mystream_b18_source_size_buf <= _mystream_b18_source_size;
        _mystream_b18_source_stride_buf <= _mystream_b18_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_52 <= _mystream_b18_source_ram_rdata;
      end 
      if((_mystream_b18_source_fsm_50 == 1) && _mystream_stream_oready) begin
        _mystream_b18_idle <= 0;
        _mystream_b18_source_ram_raddr <= _mystream_b18_source_offset_buf;
        _mystream_b18_source_ram_renable <= 1;
        _mystream_b18_source_count <= _mystream_b18_source_size_buf;
      end 
      if((_mystream_b18_source_fsm_50 == 2) && _mystream_stream_oready) begin
        _mystream_b18_source_ram_raddr <= _mystream_b18_source_ram_raddr + _mystream_b18_source_stride_buf;
        _mystream_b18_source_ram_renable <= 1;
        _mystream_b18_source_count <= _mystream_b18_source_count - 1;
      end 
      if((_mystream_b18_source_fsm_50 == 2) && (_mystream_b18_source_count == 1) && _mystream_stream_oready) begin
        _mystream_b18_source_ram_renable <= 0;
        _mystream_b18_idle <= 1;
      end 
      if((_mystream_b18_source_fsm_50 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_b18_source_ram_renable <= 0;
        _mystream_b18_idle <= 1;
      end 
      if(_set_flag_338) begin
        _mystream_b19_source_mode <= 5'b1;
        _mystream_b19_source_offset <= _th_comp_offset_4;
        _mystream_b19_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_b19_source_stride <= 1;
      end 
      if(_set_flag_338) begin
        _mystream_b19_source_sel <= 52;
      end 
      if(_mystream_source_start && _mystream_b19_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_b19_source_offset_buf <= _mystream_b19_source_offset;
        _mystream_b19_source_size_buf <= _mystream_b19_source_size;
        _mystream_b19_source_stride_buf <= _mystream_b19_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_53 <= _mystream_b19_source_ram_rdata;
      end 
      if((_mystream_b19_source_fsm_51 == 1) && _mystream_stream_oready) begin
        _mystream_b19_idle <= 0;
        _mystream_b19_source_ram_raddr <= _mystream_b19_source_offset_buf;
        _mystream_b19_source_ram_renable <= 1;
        _mystream_b19_source_count <= _mystream_b19_source_size_buf;
      end 
      if((_mystream_b19_source_fsm_51 == 2) && _mystream_stream_oready) begin
        _mystream_b19_source_ram_raddr <= _mystream_b19_source_ram_raddr + _mystream_b19_source_stride_buf;
        _mystream_b19_source_ram_renable <= 1;
        _mystream_b19_source_count <= _mystream_b19_source_count - 1;
      end 
      if((_mystream_b19_source_fsm_51 == 2) && (_mystream_b19_source_count == 1) && _mystream_stream_oready) begin
        _mystream_b19_source_ram_renable <= 0;
        _mystream_b19_idle <= 1;
      end 
      if((_mystream_b19_source_fsm_51 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_b19_source_ram_renable <= 0;
        _mystream_b19_idle <= 1;
      end 
      if(_set_flag_341) begin
        _mystream_b20_source_mode <= 5'b1;
        _mystream_b20_source_offset <= _th_comp_offset_4;
        _mystream_b20_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_b20_source_stride <= 1;
      end 
      if(_set_flag_341) begin
        _mystream_b20_source_sel <= 53;
      end 
      if(_mystream_source_start && _mystream_b20_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_b20_source_offset_buf <= _mystream_b20_source_offset;
        _mystream_b20_source_size_buf <= _mystream_b20_source_size;
        _mystream_b20_source_stride_buf <= _mystream_b20_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_54 <= _mystream_b20_source_ram_rdata;
      end 
      if((_mystream_b20_source_fsm_52 == 1) && _mystream_stream_oready) begin
        _mystream_b20_idle <= 0;
        _mystream_b20_source_ram_raddr <= _mystream_b20_source_offset_buf;
        _mystream_b20_source_ram_renable <= 1;
        _mystream_b20_source_count <= _mystream_b20_source_size_buf;
      end 
      if((_mystream_b20_source_fsm_52 == 2) && _mystream_stream_oready) begin
        _mystream_b20_source_ram_raddr <= _mystream_b20_source_ram_raddr + _mystream_b20_source_stride_buf;
        _mystream_b20_source_ram_renable <= 1;
        _mystream_b20_source_count <= _mystream_b20_source_count - 1;
      end 
      if((_mystream_b20_source_fsm_52 == 2) && (_mystream_b20_source_count == 1) && _mystream_stream_oready) begin
        _mystream_b20_source_ram_renable <= 0;
        _mystream_b20_idle <= 1;
      end 
      if((_mystream_b20_source_fsm_52 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_b20_source_ram_renable <= 0;
        _mystream_b20_idle <= 1;
      end 
      if(_set_flag_344) begin
        _mystream_b21_source_mode <= 5'b1;
        _mystream_b21_source_offset <= _th_comp_offset_4;
        _mystream_b21_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_b21_source_stride <= 1;
      end 
      if(_set_flag_344) begin
        _mystream_b21_source_sel <= 54;
      end 
      if(_mystream_source_start && _mystream_b21_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_b21_source_offset_buf <= _mystream_b21_source_offset;
        _mystream_b21_source_size_buf <= _mystream_b21_source_size;
        _mystream_b21_source_stride_buf <= _mystream_b21_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_55 <= _mystream_b21_source_ram_rdata;
      end 
      if((_mystream_b21_source_fsm_53 == 1) && _mystream_stream_oready) begin
        _mystream_b21_idle <= 0;
        _mystream_b21_source_ram_raddr <= _mystream_b21_source_offset_buf;
        _mystream_b21_source_ram_renable <= 1;
        _mystream_b21_source_count <= _mystream_b21_source_size_buf;
      end 
      if((_mystream_b21_source_fsm_53 == 2) && _mystream_stream_oready) begin
        _mystream_b21_source_ram_raddr <= _mystream_b21_source_ram_raddr + _mystream_b21_source_stride_buf;
        _mystream_b21_source_ram_renable <= 1;
        _mystream_b21_source_count <= _mystream_b21_source_count - 1;
      end 
      if((_mystream_b21_source_fsm_53 == 2) && (_mystream_b21_source_count == 1) && _mystream_stream_oready) begin
        _mystream_b21_source_ram_renable <= 0;
        _mystream_b21_idle <= 1;
      end 
      if((_mystream_b21_source_fsm_53 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_b21_source_ram_renable <= 0;
        _mystream_b21_idle <= 1;
      end 
      if(_set_flag_347) begin
        _mystream_b22_source_mode <= 5'b1;
        _mystream_b22_source_offset <= _th_comp_offset_4;
        _mystream_b22_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_b22_source_stride <= 1;
      end 
      if(_set_flag_347) begin
        _mystream_b22_source_sel <= 55;
      end 
      if(_mystream_source_start && _mystream_b22_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_b22_source_offset_buf <= _mystream_b22_source_offset;
        _mystream_b22_source_size_buf <= _mystream_b22_source_size;
        _mystream_b22_source_stride_buf <= _mystream_b22_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_56 <= _mystream_b22_source_ram_rdata;
      end 
      if((_mystream_b22_source_fsm_54 == 1) && _mystream_stream_oready) begin
        _mystream_b22_idle <= 0;
        _mystream_b22_source_ram_raddr <= _mystream_b22_source_offset_buf;
        _mystream_b22_source_ram_renable <= 1;
        _mystream_b22_source_count <= _mystream_b22_source_size_buf;
      end 
      if((_mystream_b22_source_fsm_54 == 2) && _mystream_stream_oready) begin
        _mystream_b22_source_ram_raddr <= _mystream_b22_source_ram_raddr + _mystream_b22_source_stride_buf;
        _mystream_b22_source_ram_renable <= 1;
        _mystream_b22_source_count <= _mystream_b22_source_count - 1;
      end 
      if((_mystream_b22_source_fsm_54 == 2) && (_mystream_b22_source_count == 1) && _mystream_stream_oready) begin
        _mystream_b22_source_ram_renable <= 0;
        _mystream_b22_idle <= 1;
      end 
      if((_mystream_b22_source_fsm_54 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_b22_source_ram_renable <= 0;
        _mystream_b22_idle <= 1;
      end 
      if(_set_flag_350) begin
        _mystream_b23_source_mode <= 5'b1;
        _mystream_b23_source_offset <= _th_comp_offset_4;
        _mystream_b23_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_b23_source_stride <= 1;
      end 
      if(_set_flag_350) begin
        _mystream_b23_source_sel <= 56;
      end 
      if(_mystream_source_start && _mystream_b23_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_b23_source_offset_buf <= _mystream_b23_source_offset;
        _mystream_b23_source_size_buf <= _mystream_b23_source_size;
        _mystream_b23_source_stride_buf <= _mystream_b23_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_57 <= _mystream_b23_source_ram_rdata;
      end 
      if((_mystream_b23_source_fsm_55 == 1) && _mystream_stream_oready) begin
        _mystream_b23_idle <= 0;
        _mystream_b23_source_ram_raddr <= _mystream_b23_source_offset_buf;
        _mystream_b23_source_ram_renable <= 1;
        _mystream_b23_source_count <= _mystream_b23_source_size_buf;
      end 
      if((_mystream_b23_source_fsm_55 == 2) && _mystream_stream_oready) begin
        _mystream_b23_source_ram_raddr <= _mystream_b23_source_ram_raddr + _mystream_b23_source_stride_buf;
        _mystream_b23_source_ram_renable <= 1;
        _mystream_b23_source_count <= _mystream_b23_source_count - 1;
      end 
      if((_mystream_b23_source_fsm_55 == 2) && (_mystream_b23_source_count == 1) && _mystream_stream_oready) begin
        _mystream_b23_source_ram_renable <= 0;
        _mystream_b23_idle <= 1;
      end 
      if((_mystream_b23_source_fsm_55 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_b23_source_ram_renable <= 0;
        _mystream_b23_idle <= 1;
      end 
      if(_set_flag_353) begin
        _mystream_b24_source_mode <= 5'b1;
        _mystream_b24_source_offset <= _th_comp_offset_4;
        _mystream_b24_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_b24_source_stride <= 1;
      end 
      if(_set_flag_353) begin
        _mystream_b24_source_sel <= 57;
      end 
      if(_mystream_source_start && _mystream_b24_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_b24_source_offset_buf <= _mystream_b24_source_offset;
        _mystream_b24_source_size_buf <= _mystream_b24_source_size;
        _mystream_b24_source_stride_buf <= _mystream_b24_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_58 <= _mystream_b24_source_ram_rdata;
      end 
      if((_mystream_b24_source_fsm_56 == 1) && _mystream_stream_oready) begin
        _mystream_b24_idle <= 0;
        _mystream_b24_source_ram_raddr <= _mystream_b24_source_offset_buf;
        _mystream_b24_source_ram_renable <= 1;
        _mystream_b24_source_count <= _mystream_b24_source_size_buf;
      end 
      if((_mystream_b24_source_fsm_56 == 2) && _mystream_stream_oready) begin
        _mystream_b24_source_ram_raddr <= _mystream_b24_source_ram_raddr + _mystream_b24_source_stride_buf;
        _mystream_b24_source_ram_renable <= 1;
        _mystream_b24_source_count <= _mystream_b24_source_count - 1;
      end 
      if((_mystream_b24_source_fsm_56 == 2) && (_mystream_b24_source_count == 1) && _mystream_stream_oready) begin
        _mystream_b24_source_ram_renable <= 0;
        _mystream_b24_idle <= 1;
      end 
      if((_mystream_b24_source_fsm_56 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_b24_source_ram_renable <= 0;
        _mystream_b24_idle <= 1;
      end 
      if(_set_flag_356) begin
        _mystream_b25_source_mode <= 5'b1;
        _mystream_b25_source_offset <= _th_comp_offset_4;
        _mystream_b25_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_b25_source_stride <= 1;
      end 
      if(_set_flag_356) begin
        _mystream_b25_source_sel <= 58;
      end 
      if(_mystream_source_start && _mystream_b25_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_b25_source_offset_buf <= _mystream_b25_source_offset;
        _mystream_b25_source_size_buf <= _mystream_b25_source_size;
        _mystream_b25_source_stride_buf <= _mystream_b25_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_59 <= _mystream_b25_source_ram_rdata;
      end 
      if((_mystream_b25_source_fsm_57 == 1) && _mystream_stream_oready) begin
        _mystream_b25_idle <= 0;
        _mystream_b25_source_ram_raddr <= _mystream_b25_source_offset_buf;
        _mystream_b25_source_ram_renable <= 1;
        _mystream_b25_source_count <= _mystream_b25_source_size_buf;
      end 
      if((_mystream_b25_source_fsm_57 == 2) && _mystream_stream_oready) begin
        _mystream_b25_source_ram_raddr <= _mystream_b25_source_ram_raddr + _mystream_b25_source_stride_buf;
        _mystream_b25_source_ram_renable <= 1;
        _mystream_b25_source_count <= _mystream_b25_source_count - 1;
      end 
      if((_mystream_b25_source_fsm_57 == 2) && (_mystream_b25_source_count == 1) && _mystream_stream_oready) begin
        _mystream_b25_source_ram_renable <= 0;
        _mystream_b25_idle <= 1;
      end 
      if((_mystream_b25_source_fsm_57 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_b25_source_ram_renable <= 0;
        _mystream_b25_idle <= 1;
      end 
      if(_set_flag_359) begin
        _mystream_b26_source_mode <= 5'b1;
        _mystream_b26_source_offset <= _th_comp_offset_4;
        _mystream_b26_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_b26_source_stride <= 1;
      end 
      if(_set_flag_359) begin
        _mystream_b26_source_sel <= 59;
      end 
      if(_mystream_source_start && _mystream_b26_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_b26_source_offset_buf <= _mystream_b26_source_offset;
        _mystream_b26_source_size_buf <= _mystream_b26_source_size;
        _mystream_b26_source_stride_buf <= _mystream_b26_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_60 <= _mystream_b26_source_ram_rdata;
      end 
      if((_mystream_b26_source_fsm_58 == 1) && _mystream_stream_oready) begin
        _mystream_b26_idle <= 0;
        _mystream_b26_source_ram_raddr <= _mystream_b26_source_offset_buf;
        _mystream_b26_source_ram_renable <= 1;
        _mystream_b26_source_count <= _mystream_b26_source_size_buf;
      end 
      if((_mystream_b26_source_fsm_58 == 2) && _mystream_stream_oready) begin
        _mystream_b26_source_ram_raddr <= _mystream_b26_source_ram_raddr + _mystream_b26_source_stride_buf;
        _mystream_b26_source_ram_renable <= 1;
        _mystream_b26_source_count <= _mystream_b26_source_count - 1;
      end 
      if((_mystream_b26_source_fsm_58 == 2) && (_mystream_b26_source_count == 1) && _mystream_stream_oready) begin
        _mystream_b26_source_ram_renable <= 0;
        _mystream_b26_idle <= 1;
      end 
      if((_mystream_b26_source_fsm_58 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_b26_source_ram_renable <= 0;
        _mystream_b26_idle <= 1;
      end 
      if(_set_flag_362) begin
        _mystream_b27_source_mode <= 5'b1;
        _mystream_b27_source_offset <= _th_comp_offset_4;
        _mystream_b27_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_b27_source_stride <= 1;
      end 
      if(_set_flag_362) begin
        _mystream_b27_source_sel <= 60;
      end 
      if(_mystream_source_start && _mystream_b27_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_b27_source_offset_buf <= _mystream_b27_source_offset;
        _mystream_b27_source_size_buf <= _mystream_b27_source_size;
        _mystream_b27_source_stride_buf <= _mystream_b27_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_61 <= _mystream_b27_source_ram_rdata;
      end 
      if((_mystream_b27_source_fsm_59 == 1) && _mystream_stream_oready) begin
        _mystream_b27_idle <= 0;
        _mystream_b27_source_ram_raddr <= _mystream_b27_source_offset_buf;
        _mystream_b27_source_ram_renable <= 1;
        _mystream_b27_source_count <= _mystream_b27_source_size_buf;
      end 
      if((_mystream_b27_source_fsm_59 == 2) && _mystream_stream_oready) begin
        _mystream_b27_source_ram_raddr <= _mystream_b27_source_ram_raddr + _mystream_b27_source_stride_buf;
        _mystream_b27_source_ram_renable <= 1;
        _mystream_b27_source_count <= _mystream_b27_source_count - 1;
      end 
      if((_mystream_b27_source_fsm_59 == 2) && (_mystream_b27_source_count == 1) && _mystream_stream_oready) begin
        _mystream_b27_source_ram_renable <= 0;
        _mystream_b27_idle <= 1;
      end 
      if((_mystream_b27_source_fsm_59 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_b27_source_ram_renable <= 0;
        _mystream_b27_idle <= 1;
      end 
      if(_set_flag_365) begin
        _mystream_b28_source_mode <= 5'b1;
        _mystream_b28_source_offset <= _th_comp_offset_4;
        _mystream_b28_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_b28_source_stride <= 1;
      end 
      if(_set_flag_365) begin
        _mystream_b28_source_sel <= 61;
      end 
      if(_mystream_source_start && _mystream_b28_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_b28_source_offset_buf <= _mystream_b28_source_offset;
        _mystream_b28_source_size_buf <= _mystream_b28_source_size;
        _mystream_b28_source_stride_buf <= _mystream_b28_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_62 <= _mystream_b28_source_ram_rdata;
      end 
      if((_mystream_b28_source_fsm_60 == 1) && _mystream_stream_oready) begin
        _mystream_b28_idle <= 0;
        _mystream_b28_source_ram_raddr <= _mystream_b28_source_offset_buf;
        _mystream_b28_source_ram_renable <= 1;
        _mystream_b28_source_count <= _mystream_b28_source_size_buf;
      end 
      if((_mystream_b28_source_fsm_60 == 2) && _mystream_stream_oready) begin
        _mystream_b28_source_ram_raddr <= _mystream_b28_source_ram_raddr + _mystream_b28_source_stride_buf;
        _mystream_b28_source_ram_renable <= 1;
        _mystream_b28_source_count <= _mystream_b28_source_count - 1;
      end 
      if((_mystream_b28_source_fsm_60 == 2) && (_mystream_b28_source_count == 1) && _mystream_stream_oready) begin
        _mystream_b28_source_ram_renable <= 0;
        _mystream_b28_idle <= 1;
      end 
      if((_mystream_b28_source_fsm_60 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_b28_source_ram_renable <= 0;
        _mystream_b28_idle <= 1;
      end 
      if(_set_flag_368) begin
        _mystream_b29_source_mode <= 5'b1;
        _mystream_b29_source_offset <= _th_comp_offset_4;
        _mystream_b29_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_b29_source_stride <= 1;
      end 
      if(_set_flag_368) begin
        _mystream_b29_source_sel <= 62;
      end 
      if(_mystream_source_start && _mystream_b29_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_b29_source_offset_buf <= _mystream_b29_source_offset;
        _mystream_b29_source_size_buf <= _mystream_b29_source_size;
        _mystream_b29_source_stride_buf <= _mystream_b29_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_63 <= _mystream_b29_source_ram_rdata;
      end 
      if((_mystream_b29_source_fsm_61 == 1) && _mystream_stream_oready) begin
        _mystream_b29_idle <= 0;
        _mystream_b29_source_ram_raddr <= _mystream_b29_source_offset_buf;
        _mystream_b29_source_ram_renable <= 1;
        _mystream_b29_source_count <= _mystream_b29_source_size_buf;
      end 
      if((_mystream_b29_source_fsm_61 == 2) && _mystream_stream_oready) begin
        _mystream_b29_source_ram_raddr <= _mystream_b29_source_ram_raddr + _mystream_b29_source_stride_buf;
        _mystream_b29_source_ram_renable <= 1;
        _mystream_b29_source_count <= _mystream_b29_source_count - 1;
      end 
      if((_mystream_b29_source_fsm_61 == 2) && (_mystream_b29_source_count == 1) && _mystream_stream_oready) begin
        _mystream_b29_source_ram_renable <= 0;
        _mystream_b29_idle <= 1;
      end 
      if((_mystream_b29_source_fsm_61 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_b29_source_ram_renable <= 0;
        _mystream_b29_idle <= 1;
      end 
      if(_set_flag_371) begin
        _mystream_b30_source_mode <= 5'b1;
        _mystream_b30_source_offset <= _th_comp_offset_4;
        _mystream_b30_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_b30_source_stride <= 1;
      end 
      if(_set_flag_371) begin
        _mystream_b30_source_sel <= 63;
      end 
      if(_mystream_source_start && _mystream_b30_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_b30_source_offset_buf <= _mystream_b30_source_offset;
        _mystream_b30_source_size_buf <= _mystream_b30_source_size;
        _mystream_b30_source_stride_buf <= _mystream_b30_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_64 <= _mystream_b30_source_ram_rdata;
      end 
      if((_mystream_b30_source_fsm_62 == 1) && _mystream_stream_oready) begin
        _mystream_b30_idle <= 0;
        _mystream_b30_source_ram_raddr <= _mystream_b30_source_offset_buf;
        _mystream_b30_source_ram_renable <= 1;
        _mystream_b30_source_count <= _mystream_b30_source_size_buf;
      end 
      if((_mystream_b30_source_fsm_62 == 2) && _mystream_stream_oready) begin
        _mystream_b30_source_ram_raddr <= _mystream_b30_source_ram_raddr + _mystream_b30_source_stride_buf;
        _mystream_b30_source_ram_renable <= 1;
        _mystream_b30_source_count <= _mystream_b30_source_count - 1;
      end 
      if((_mystream_b30_source_fsm_62 == 2) && (_mystream_b30_source_count == 1) && _mystream_stream_oready) begin
        _mystream_b30_source_ram_renable <= 0;
        _mystream_b30_idle <= 1;
      end 
      if((_mystream_b30_source_fsm_62 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_b30_source_ram_renable <= 0;
        _mystream_b30_idle <= 1;
      end 
      if(_set_flag_374) begin
        _mystream_b31_source_mode <= 5'b1;
        _mystream_b31_source_offset <= _th_comp_offset_4;
        _mystream_b31_source_size <= _th_comp_size_3 + 32 - 1 >>> 5;
        _mystream_b31_source_stride <= 1;
      end 
      if(_set_flag_374) begin
        _mystream_b31_source_sel <= 64;
      end 
      if(_mystream_source_start && _mystream_b31_source_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_b31_source_offset_buf <= _mystream_b31_source_offset;
        _mystream_b31_source_size_buf <= _mystream_b31_source_size;
        _mystream_b31_source_stride_buf <= _mystream_b31_source_stride;
      end 
      if(_mystream_stream_oready && _mystream_source_busy && _mystream_is_root) begin
        __variable_wdata_65 <= _mystream_b31_source_ram_rdata;
      end 
      if((_mystream_b31_source_fsm_63 == 1) && _mystream_stream_oready) begin
        _mystream_b31_idle <= 0;
        _mystream_b31_source_ram_raddr <= _mystream_b31_source_offset_buf;
        _mystream_b31_source_ram_renable <= 1;
        _mystream_b31_source_count <= _mystream_b31_source_size_buf;
      end 
      if((_mystream_b31_source_fsm_63 == 2) && _mystream_stream_oready) begin
        _mystream_b31_source_ram_raddr <= _mystream_b31_source_ram_raddr + _mystream_b31_source_stride_buf;
        _mystream_b31_source_ram_renable <= 1;
        _mystream_b31_source_count <= _mystream_b31_source_count - 1;
      end 
      if((_mystream_b31_source_fsm_63 == 2) && (_mystream_b31_source_count == 1) && _mystream_stream_oready) begin
        _mystream_b31_source_ram_renable <= 0;
        _mystream_b31_idle <= 1;
      end 
      if((_mystream_b31_source_fsm_63 == 2) && _mystream_source_stop && _mystream_stream_oready) begin
        _mystream_b31_source_ram_renable <= 0;
        _mystream_b31_idle <= 1;
      end 
      if(_mystream_stream_oready) begin
        _tmp_378 <= _set_flag_377;
      end 
      if(_mystream_stream_oready) begin
        _tmp_379 <= _tmp_378;
      end 
      if(_mystream_stream_oready) begin
        _tmp_380 <= _tmp_379;
      end 
      if(_mystream_stream_oready) begin
        _tmp_381 <= _tmp_380;
      end 
      if(_mystream_stream_oready) begin
        _tmp_382 <= _tmp_381;
      end 
      if(_mystream_stream_oready) begin
        _tmp_383 <= _tmp_382;
      end 
      if(_mystream_stream_oready) begin
        _tmp_384 <= _th_comp_offset_4;
      end 
      if(_mystream_stream_oready) begin
        _tmp_385 <= _tmp_384;
      end 
      if(_mystream_stream_oready) begin
        _tmp_386 <= _tmp_385;
      end 
      if(_mystream_stream_oready) begin
        _tmp_387 <= _tmp_386;
      end 
      if(_mystream_stream_oready) begin
        _tmp_388 <= _tmp_387;
      end 
      if(_mystream_stream_oready) begin
        _tmp_389 <= _tmp_388;
      end 
      if(_mystream_stream_oready) begin
        _tmp_392 <= _tmp_391;
      end 
      if(_mystream_stream_oready) begin
        _tmp_393 <= _tmp_392;
      end 
      if(_mystream_stream_oready) begin
        _tmp_394 <= _tmp_393;
      end 
      if(_mystream_stream_oready) begin
        _tmp_395 <= _tmp_394;
      end 
      if(_mystream_stream_oready) begin
        _tmp_396 <= _tmp_395;
      end 
      if(_mystream_stream_oready) begin
        _tmp_397 <= _tmp_396;
      end 
      if(_tmp_383) begin
        _mystream_sum_vec0_sink_mode <= 5'b1;
        _mystream_sum_vec0_sink_offset <= _tmp_389;
        _mystream_sum_vec0_sink_size <= _tmp_397;
        _mystream_sum_vec0_sink_stride <= 1;
      end 
      if(_tmp_383) begin
        _mystream_sum_vec0_sink_sel <= 65;
      end 
      if(_mystream_sink_start && _mystream_sum_vec0_sink_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_sum_vec0_sink_offset_buf <= _mystream_sum_vec0_sink_offset;
        _mystream_sum_vec0_sink_size_buf <= _mystream_sum_vec0_sink_size;
        _mystream_sum_vec0_sink_stride_buf <= _mystream_sum_vec0_sink_stride;
      end 
      if((_mystream_sum_vec0_sink_fsm_64 == 1) && _mystream_stream_oready) begin
        _mystream_sum_vec0_sink_waddr <= _mystream_sum_vec0_sink_offset_buf - _mystream_sum_vec0_sink_stride_buf;
        _mystream_sum_vec0_sink_count <= _mystream_sum_vec0_sink_size_buf;
      end 
      if((_mystream_sum_vec0_sink_fsm_64 == 2) && _mystream_stream_oready) begin
        _mystream_sum_vec0_sink_waddr <= _mystream_sum_vec0_sink_waddr + _mystream_sum_vec0_sink_stride_buf;
        _mystream_sum_vec0_sink_wdata <= mystream_sum_vec0_data;
        _mystream_sum_vec0_sink_wenable <= 1;
        _mystream_sum_vec0_sink_count <= _mystream_sum_vec0_sink_count - 1;
      end 
      if(_mystream_stream_oready) begin
        _tmp_399 <= _set_flag_398;
      end 
      if(_mystream_stream_oready) begin
        _tmp_400 <= _tmp_399;
      end 
      if(_mystream_stream_oready) begin
        _tmp_401 <= _tmp_400;
      end 
      if(_mystream_stream_oready) begin
        _tmp_402 <= _tmp_401;
      end 
      if(_mystream_stream_oready) begin
        _tmp_403 <= _tmp_402;
      end 
      if(_mystream_stream_oready) begin
        _tmp_404 <= _tmp_403;
      end 
      if(_mystream_stream_oready) begin
        _tmp_405 <= _th_comp_offset_4;
      end 
      if(_mystream_stream_oready) begin
        _tmp_406 <= _tmp_405;
      end 
      if(_mystream_stream_oready) begin
        _tmp_407 <= _tmp_406;
      end 
      if(_mystream_stream_oready) begin
        _tmp_408 <= _tmp_407;
      end 
      if(_mystream_stream_oready) begin
        _tmp_409 <= _tmp_408;
      end 
      if(_mystream_stream_oready) begin
        _tmp_410 <= _tmp_409;
      end 
      if(_mystream_stream_oready) begin
        _tmp_413 <= _tmp_412;
      end 
      if(_mystream_stream_oready) begin
        _tmp_414 <= _tmp_413;
      end 
      if(_mystream_stream_oready) begin
        _tmp_415 <= _tmp_414;
      end 
      if(_mystream_stream_oready) begin
        _tmp_416 <= _tmp_415;
      end 
      if(_mystream_stream_oready) begin
        _tmp_417 <= _tmp_416;
      end 
      if(_mystream_stream_oready) begin
        _tmp_418 <= _tmp_417;
      end 
      if(_tmp_404) begin
        _mystream_sum_vec1_sink_mode <= 5'b1;
        _mystream_sum_vec1_sink_offset <= _tmp_410;
        _mystream_sum_vec1_sink_size <= _tmp_418;
        _mystream_sum_vec1_sink_stride <= 1;
      end 
      if(_tmp_404) begin
        _mystream_sum_vec1_sink_sel <= 66;
      end 
      if(_mystream_sink_start && _mystream_sum_vec1_sink_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_sum_vec1_sink_offset_buf <= _mystream_sum_vec1_sink_offset;
        _mystream_sum_vec1_sink_size_buf <= _mystream_sum_vec1_sink_size;
        _mystream_sum_vec1_sink_stride_buf <= _mystream_sum_vec1_sink_stride;
      end 
      if((_mystream_sum_vec1_sink_fsm_65 == 1) && _mystream_stream_oready) begin
        _mystream_sum_vec1_sink_waddr <= _mystream_sum_vec1_sink_offset_buf - _mystream_sum_vec1_sink_stride_buf;
        _mystream_sum_vec1_sink_count <= _mystream_sum_vec1_sink_size_buf;
      end 
      if((_mystream_sum_vec1_sink_fsm_65 == 2) && _mystream_stream_oready) begin
        _mystream_sum_vec1_sink_waddr <= _mystream_sum_vec1_sink_waddr + _mystream_sum_vec1_sink_stride_buf;
        _mystream_sum_vec1_sink_wdata <= mystream_sum_vec1_data;
        _mystream_sum_vec1_sink_wenable <= 1;
        _mystream_sum_vec1_sink_count <= _mystream_sum_vec1_sink_count - 1;
      end 
      if(_mystream_stream_oready) begin
        _tmp_420 <= _set_flag_419;
      end 
      if(_mystream_stream_oready) begin
        _tmp_421 <= _tmp_420;
      end 
      if(_mystream_stream_oready) begin
        _tmp_422 <= _tmp_421;
      end 
      if(_mystream_stream_oready) begin
        _tmp_423 <= _tmp_422;
      end 
      if(_mystream_stream_oready) begin
        _tmp_424 <= _tmp_423;
      end 
      if(_mystream_stream_oready) begin
        _tmp_425 <= _tmp_424;
      end 
      if(_mystream_stream_oready) begin
        _tmp_426 <= _th_comp_offset_4;
      end 
      if(_mystream_stream_oready) begin
        _tmp_427 <= _tmp_426;
      end 
      if(_mystream_stream_oready) begin
        _tmp_428 <= _tmp_427;
      end 
      if(_mystream_stream_oready) begin
        _tmp_429 <= _tmp_428;
      end 
      if(_mystream_stream_oready) begin
        _tmp_430 <= _tmp_429;
      end 
      if(_mystream_stream_oready) begin
        _tmp_431 <= _tmp_430;
      end 
      if(_mystream_stream_oready) begin
        _tmp_434 <= _tmp_433;
      end 
      if(_mystream_stream_oready) begin
        _tmp_435 <= _tmp_434;
      end 
      if(_mystream_stream_oready) begin
        _tmp_436 <= _tmp_435;
      end 
      if(_mystream_stream_oready) begin
        _tmp_437 <= _tmp_436;
      end 
      if(_mystream_stream_oready) begin
        _tmp_438 <= _tmp_437;
      end 
      if(_mystream_stream_oready) begin
        _tmp_439 <= _tmp_438;
      end 
      if(_tmp_425) begin
        _mystream_sum_vec2_sink_mode <= 5'b1;
        _mystream_sum_vec2_sink_offset <= _tmp_431;
        _mystream_sum_vec2_sink_size <= _tmp_439;
        _mystream_sum_vec2_sink_stride <= 1;
      end 
      if(_tmp_425) begin
        _mystream_sum_vec2_sink_sel <= 67;
      end 
      if(_mystream_sink_start && _mystream_sum_vec2_sink_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_sum_vec2_sink_offset_buf <= _mystream_sum_vec2_sink_offset;
        _mystream_sum_vec2_sink_size_buf <= _mystream_sum_vec2_sink_size;
        _mystream_sum_vec2_sink_stride_buf <= _mystream_sum_vec2_sink_stride;
      end 
      if((_mystream_sum_vec2_sink_fsm_66 == 1) && _mystream_stream_oready) begin
        _mystream_sum_vec2_sink_waddr <= _mystream_sum_vec2_sink_offset_buf - _mystream_sum_vec2_sink_stride_buf;
        _mystream_sum_vec2_sink_count <= _mystream_sum_vec2_sink_size_buf;
      end 
      if((_mystream_sum_vec2_sink_fsm_66 == 2) && _mystream_stream_oready) begin
        _mystream_sum_vec2_sink_waddr <= _mystream_sum_vec2_sink_waddr + _mystream_sum_vec2_sink_stride_buf;
        _mystream_sum_vec2_sink_wdata <= mystream_sum_vec2_data;
        _mystream_sum_vec2_sink_wenable <= 1;
        _mystream_sum_vec2_sink_count <= _mystream_sum_vec2_sink_count - 1;
      end 
      if(_mystream_stream_oready) begin
        _tmp_441 <= _set_flag_440;
      end 
      if(_mystream_stream_oready) begin
        _tmp_442 <= _tmp_441;
      end 
      if(_mystream_stream_oready) begin
        _tmp_443 <= _tmp_442;
      end 
      if(_mystream_stream_oready) begin
        _tmp_444 <= _tmp_443;
      end 
      if(_mystream_stream_oready) begin
        _tmp_445 <= _tmp_444;
      end 
      if(_mystream_stream_oready) begin
        _tmp_446 <= _tmp_445;
      end 
      if(_mystream_stream_oready) begin
        _tmp_447 <= _th_comp_offset_4;
      end 
      if(_mystream_stream_oready) begin
        _tmp_448 <= _tmp_447;
      end 
      if(_mystream_stream_oready) begin
        _tmp_449 <= _tmp_448;
      end 
      if(_mystream_stream_oready) begin
        _tmp_450 <= _tmp_449;
      end 
      if(_mystream_stream_oready) begin
        _tmp_451 <= _tmp_450;
      end 
      if(_mystream_stream_oready) begin
        _tmp_452 <= _tmp_451;
      end 
      if(_mystream_stream_oready) begin
        _tmp_455 <= _tmp_454;
      end 
      if(_mystream_stream_oready) begin
        _tmp_456 <= _tmp_455;
      end 
      if(_mystream_stream_oready) begin
        _tmp_457 <= _tmp_456;
      end 
      if(_mystream_stream_oready) begin
        _tmp_458 <= _tmp_457;
      end 
      if(_mystream_stream_oready) begin
        _tmp_459 <= _tmp_458;
      end 
      if(_mystream_stream_oready) begin
        _tmp_460 <= _tmp_459;
      end 
      if(_tmp_446) begin
        _mystream_sum_vec3_sink_mode <= 5'b1;
        _mystream_sum_vec3_sink_offset <= _tmp_452;
        _mystream_sum_vec3_sink_size <= _tmp_460;
        _mystream_sum_vec3_sink_stride <= 1;
      end 
      if(_tmp_446) begin
        _mystream_sum_vec3_sink_sel <= 68;
      end 
      if(_mystream_sink_start && _mystream_sum_vec3_sink_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_sum_vec3_sink_offset_buf <= _mystream_sum_vec3_sink_offset;
        _mystream_sum_vec3_sink_size_buf <= _mystream_sum_vec3_sink_size;
        _mystream_sum_vec3_sink_stride_buf <= _mystream_sum_vec3_sink_stride;
      end 
      if((_mystream_sum_vec3_sink_fsm_67 == 1) && _mystream_stream_oready) begin
        _mystream_sum_vec3_sink_waddr <= _mystream_sum_vec3_sink_offset_buf - _mystream_sum_vec3_sink_stride_buf;
        _mystream_sum_vec3_sink_count <= _mystream_sum_vec3_sink_size_buf;
      end 
      if((_mystream_sum_vec3_sink_fsm_67 == 2) && _mystream_stream_oready) begin
        _mystream_sum_vec3_sink_waddr <= _mystream_sum_vec3_sink_waddr + _mystream_sum_vec3_sink_stride_buf;
        _mystream_sum_vec3_sink_wdata <= mystream_sum_vec3_data;
        _mystream_sum_vec3_sink_wenable <= 1;
        _mystream_sum_vec3_sink_count <= _mystream_sum_vec3_sink_count - 1;
      end 
      if(_mystream_stream_oready) begin
        _tmp_462 <= _set_flag_461;
      end 
      if(_mystream_stream_oready) begin
        _tmp_463 <= _tmp_462;
      end 
      if(_mystream_stream_oready) begin
        _tmp_464 <= _tmp_463;
      end 
      if(_mystream_stream_oready) begin
        _tmp_465 <= _tmp_464;
      end 
      if(_mystream_stream_oready) begin
        _tmp_466 <= _tmp_465;
      end 
      if(_mystream_stream_oready) begin
        _tmp_467 <= _tmp_466;
      end 
      if(_mystream_stream_oready) begin
        _tmp_468 <= _th_comp_offset_4;
      end 
      if(_mystream_stream_oready) begin
        _tmp_469 <= _tmp_468;
      end 
      if(_mystream_stream_oready) begin
        _tmp_470 <= _tmp_469;
      end 
      if(_mystream_stream_oready) begin
        _tmp_471 <= _tmp_470;
      end 
      if(_mystream_stream_oready) begin
        _tmp_472 <= _tmp_471;
      end 
      if(_mystream_stream_oready) begin
        _tmp_473 <= _tmp_472;
      end 
      if(_mystream_stream_oready) begin
        _tmp_476 <= _tmp_475;
      end 
      if(_mystream_stream_oready) begin
        _tmp_477 <= _tmp_476;
      end 
      if(_mystream_stream_oready) begin
        _tmp_478 <= _tmp_477;
      end 
      if(_mystream_stream_oready) begin
        _tmp_479 <= _tmp_478;
      end 
      if(_mystream_stream_oready) begin
        _tmp_480 <= _tmp_479;
      end 
      if(_mystream_stream_oready) begin
        _tmp_481 <= _tmp_480;
      end 
      if(_tmp_467) begin
        _mystream_sum_vec4_sink_mode <= 5'b1;
        _mystream_sum_vec4_sink_offset <= _tmp_473;
        _mystream_sum_vec4_sink_size <= _tmp_481;
        _mystream_sum_vec4_sink_stride <= 1;
      end 
      if(_tmp_467) begin
        _mystream_sum_vec4_sink_sel <= 69;
      end 
      if(_mystream_sink_start && _mystream_sum_vec4_sink_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_sum_vec4_sink_offset_buf <= _mystream_sum_vec4_sink_offset;
        _mystream_sum_vec4_sink_size_buf <= _mystream_sum_vec4_sink_size;
        _mystream_sum_vec4_sink_stride_buf <= _mystream_sum_vec4_sink_stride;
      end 
      if((_mystream_sum_vec4_sink_fsm_68 == 1) && _mystream_stream_oready) begin
        _mystream_sum_vec4_sink_waddr <= _mystream_sum_vec4_sink_offset_buf - _mystream_sum_vec4_sink_stride_buf;
        _mystream_sum_vec4_sink_count <= _mystream_sum_vec4_sink_size_buf;
      end 
      if((_mystream_sum_vec4_sink_fsm_68 == 2) && _mystream_stream_oready) begin
        _mystream_sum_vec4_sink_waddr <= _mystream_sum_vec4_sink_waddr + _mystream_sum_vec4_sink_stride_buf;
        _mystream_sum_vec4_sink_wdata <= mystream_sum_vec4_data;
        _mystream_sum_vec4_sink_wenable <= 1;
        _mystream_sum_vec4_sink_count <= _mystream_sum_vec4_sink_count - 1;
      end 
      if(_mystream_stream_oready) begin
        _tmp_483 <= _set_flag_482;
      end 
      if(_mystream_stream_oready) begin
        _tmp_484 <= _tmp_483;
      end 
      if(_mystream_stream_oready) begin
        _tmp_485 <= _tmp_484;
      end 
      if(_mystream_stream_oready) begin
        _tmp_486 <= _tmp_485;
      end 
      if(_mystream_stream_oready) begin
        _tmp_487 <= _tmp_486;
      end 
      if(_mystream_stream_oready) begin
        _tmp_488 <= _tmp_487;
      end 
      if(_mystream_stream_oready) begin
        _tmp_489 <= _th_comp_offset_4;
      end 
      if(_mystream_stream_oready) begin
        _tmp_490 <= _tmp_489;
      end 
      if(_mystream_stream_oready) begin
        _tmp_491 <= _tmp_490;
      end 
      if(_mystream_stream_oready) begin
        _tmp_492 <= _tmp_491;
      end 
      if(_mystream_stream_oready) begin
        _tmp_493 <= _tmp_492;
      end 
      if(_mystream_stream_oready) begin
        _tmp_494 <= _tmp_493;
      end 
      if(_mystream_stream_oready) begin
        _tmp_497 <= _tmp_496;
      end 
      if(_mystream_stream_oready) begin
        _tmp_498 <= _tmp_497;
      end 
      if(_mystream_stream_oready) begin
        _tmp_499 <= _tmp_498;
      end 
      if(_mystream_stream_oready) begin
        _tmp_500 <= _tmp_499;
      end 
      if(_mystream_stream_oready) begin
        _tmp_501 <= _tmp_500;
      end 
      if(_mystream_stream_oready) begin
        _tmp_502 <= _tmp_501;
      end 
      if(_tmp_488) begin
        _mystream_sum_vec5_sink_mode <= 5'b1;
        _mystream_sum_vec5_sink_offset <= _tmp_494;
        _mystream_sum_vec5_sink_size <= _tmp_502;
        _mystream_sum_vec5_sink_stride <= 1;
      end 
      if(_tmp_488) begin
        _mystream_sum_vec5_sink_sel <= 70;
      end 
      if(_mystream_sink_start && _mystream_sum_vec5_sink_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_sum_vec5_sink_offset_buf <= _mystream_sum_vec5_sink_offset;
        _mystream_sum_vec5_sink_size_buf <= _mystream_sum_vec5_sink_size;
        _mystream_sum_vec5_sink_stride_buf <= _mystream_sum_vec5_sink_stride;
      end 
      if((_mystream_sum_vec5_sink_fsm_69 == 1) && _mystream_stream_oready) begin
        _mystream_sum_vec5_sink_waddr <= _mystream_sum_vec5_sink_offset_buf - _mystream_sum_vec5_sink_stride_buf;
        _mystream_sum_vec5_sink_count <= _mystream_sum_vec5_sink_size_buf;
      end 
      if((_mystream_sum_vec5_sink_fsm_69 == 2) && _mystream_stream_oready) begin
        _mystream_sum_vec5_sink_waddr <= _mystream_sum_vec5_sink_waddr + _mystream_sum_vec5_sink_stride_buf;
        _mystream_sum_vec5_sink_wdata <= mystream_sum_vec5_data;
        _mystream_sum_vec5_sink_wenable <= 1;
        _mystream_sum_vec5_sink_count <= _mystream_sum_vec5_sink_count - 1;
      end 
      if(_mystream_stream_oready) begin
        _tmp_504 <= _set_flag_503;
      end 
      if(_mystream_stream_oready) begin
        _tmp_505 <= _tmp_504;
      end 
      if(_mystream_stream_oready) begin
        _tmp_506 <= _tmp_505;
      end 
      if(_mystream_stream_oready) begin
        _tmp_507 <= _tmp_506;
      end 
      if(_mystream_stream_oready) begin
        _tmp_508 <= _tmp_507;
      end 
      if(_mystream_stream_oready) begin
        _tmp_509 <= _tmp_508;
      end 
      if(_mystream_stream_oready) begin
        _tmp_510 <= _th_comp_offset_4;
      end 
      if(_mystream_stream_oready) begin
        _tmp_511 <= _tmp_510;
      end 
      if(_mystream_stream_oready) begin
        _tmp_512 <= _tmp_511;
      end 
      if(_mystream_stream_oready) begin
        _tmp_513 <= _tmp_512;
      end 
      if(_mystream_stream_oready) begin
        _tmp_514 <= _tmp_513;
      end 
      if(_mystream_stream_oready) begin
        _tmp_515 <= _tmp_514;
      end 
      if(_mystream_stream_oready) begin
        _tmp_518 <= _tmp_517;
      end 
      if(_mystream_stream_oready) begin
        _tmp_519 <= _tmp_518;
      end 
      if(_mystream_stream_oready) begin
        _tmp_520 <= _tmp_519;
      end 
      if(_mystream_stream_oready) begin
        _tmp_521 <= _tmp_520;
      end 
      if(_mystream_stream_oready) begin
        _tmp_522 <= _tmp_521;
      end 
      if(_mystream_stream_oready) begin
        _tmp_523 <= _tmp_522;
      end 
      if(_tmp_509) begin
        _mystream_sum_vec6_sink_mode <= 5'b1;
        _mystream_sum_vec6_sink_offset <= _tmp_515;
        _mystream_sum_vec6_sink_size <= _tmp_523;
        _mystream_sum_vec6_sink_stride <= 1;
      end 
      if(_tmp_509) begin
        _mystream_sum_vec6_sink_sel <= 71;
      end 
      if(_mystream_sink_start && _mystream_sum_vec6_sink_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_sum_vec6_sink_offset_buf <= _mystream_sum_vec6_sink_offset;
        _mystream_sum_vec6_sink_size_buf <= _mystream_sum_vec6_sink_size;
        _mystream_sum_vec6_sink_stride_buf <= _mystream_sum_vec6_sink_stride;
      end 
      if((_mystream_sum_vec6_sink_fsm_70 == 1) && _mystream_stream_oready) begin
        _mystream_sum_vec6_sink_waddr <= _mystream_sum_vec6_sink_offset_buf - _mystream_sum_vec6_sink_stride_buf;
        _mystream_sum_vec6_sink_count <= _mystream_sum_vec6_sink_size_buf;
      end 
      if((_mystream_sum_vec6_sink_fsm_70 == 2) && _mystream_stream_oready) begin
        _mystream_sum_vec6_sink_waddr <= _mystream_sum_vec6_sink_waddr + _mystream_sum_vec6_sink_stride_buf;
        _mystream_sum_vec6_sink_wdata <= mystream_sum_vec6_data;
        _mystream_sum_vec6_sink_wenable <= 1;
        _mystream_sum_vec6_sink_count <= _mystream_sum_vec6_sink_count - 1;
      end 
      if(_mystream_stream_oready) begin
        _tmp_525 <= _set_flag_524;
      end 
      if(_mystream_stream_oready) begin
        _tmp_526 <= _tmp_525;
      end 
      if(_mystream_stream_oready) begin
        _tmp_527 <= _tmp_526;
      end 
      if(_mystream_stream_oready) begin
        _tmp_528 <= _tmp_527;
      end 
      if(_mystream_stream_oready) begin
        _tmp_529 <= _tmp_528;
      end 
      if(_mystream_stream_oready) begin
        _tmp_530 <= _tmp_529;
      end 
      if(_mystream_stream_oready) begin
        _tmp_531 <= _th_comp_offset_4;
      end 
      if(_mystream_stream_oready) begin
        _tmp_532 <= _tmp_531;
      end 
      if(_mystream_stream_oready) begin
        _tmp_533 <= _tmp_532;
      end 
      if(_mystream_stream_oready) begin
        _tmp_534 <= _tmp_533;
      end 
      if(_mystream_stream_oready) begin
        _tmp_535 <= _tmp_534;
      end 
      if(_mystream_stream_oready) begin
        _tmp_536 <= _tmp_535;
      end 
      if(_mystream_stream_oready) begin
        _tmp_539 <= _tmp_538;
      end 
      if(_mystream_stream_oready) begin
        _tmp_540 <= _tmp_539;
      end 
      if(_mystream_stream_oready) begin
        _tmp_541 <= _tmp_540;
      end 
      if(_mystream_stream_oready) begin
        _tmp_542 <= _tmp_541;
      end 
      if(_mystream_stream_oready) begin
        _tmp_543 <= _tmp_542;
      end 
      if(_mystream_stream_oready) begin
        _tmp_544 <= _tmp_543;
      end 
      if(_tmp_530) begin
        _mystream_sum_vec7_sink_mode <= 5'b1;
        _mystream_sum_vec7_sink_offset <= _tmp_536;
        _mystream_sum_vec7_sink_size <= _tmp_544;
        _mystream_sum_vec7_sink_stride <= 1;
      end 
      if(_tmp_530) begin
        _mystream_sum_vec7_sink_sel <= 72;
      end 
      if(_mystream_sink_start && _mystream_sum_vec7_sink_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_sum_vec7_sink_offset_buf <= _mystream_sum_vec7_sink_offset;
        _mystream_sum_vec7_sink_size_buf <= _mystream_sum_vec7_sink_size;
        _mystream_sum_vec7_sink_stride_buf <= _mystream_sum_vec7_sink_stride;
      end 
      if((_mystream_sum_vec7_sink_fsm_71 == 1) && _mystream_stream_oready) begin
        _mystream_sum_vec7_sink_waddr <= _mystream_sum_vec7_sink_offset_buf - _mystream_sum_vec7_sink_stride_buf;
        _mystream_sum_vec7_sink_count <= _mystream_sum_vec7_sink_size_buf;
      end 
      if((_mystream_sum_vec7_sink_fsm_71 == 2) && _mystream_stream_oready) begin
        _mystream_sum_vec7_sink_waddr <= _mystream_sum_vec7_sink_waddr + _mystream_sum_vec7_sink_stride_buf;
        _mystream_sum_vec7_sink_wdata <= mystream_sum_vec7_data;
        _mystream_sum_vec7_sink_wenable <= 1;
        _mystream_sum_vec7_sink_count <= _mystream_sum_vec7_sink_count - 1;
      end 
      if(_mystream_stream_oready) begin
        _tmp_546 <= _set_flag_545;
      end 
      if(_mystream_stream_oready) begin
        _tmp_547 <= _tmp_546;
      end 
      if(_mystream_stream_oready) begin
        _tmp_548 <= _tmp_547;
      end 
      if(_mystream_stream_oready) begin
        _tmp_549 <= _tmp_548;
      end 
      if(_mystream_stream_oready) begin
        _tmp_550 <= _tmp_549;
      end 
      if(_mystream_stream_oready) begin
        _tmp_551 <= _tmp_550;
      end 
      if(_mystream_stream_oready) begin
        _tmp_552 <= _th_comp_offset_4;
      end 
      if(_mystream_stream_oready) begin
        _tmp_553 <= _tmp_552;
      end 
      if(_mystream_stream_oready) begin
        _tmp_554 <= _tmp_553;
      end 
      if(_mystream_stream_oready) begin
        _tmp_555 <= _tmp_554;
      end 
      if(_mystream_stream_oready) begin
        _tmp_556 <= _tmp_555;
      end 
      if(_mystream_stream_oready) begin
        _tmp_557 <= _tmp_556;
      end 
      if(_mystream_stream_oready) begin
        _tmp_560 <= _tmp_559;
      end 
      if(_mystream_stream_oready) begin
        _tmp_561 <= _tmp_560;
      end 
      if(_mystream_stream_oready) begin
        _tmp_562 <= _tmp_561;
      end 
      if(_mystream_stream_oready) begin
        _tmp_563 <= _tmp_562;
      end 
      if(_mystream_stream_oready) begin
        _tmp_564 <= _tmp_563;
      end 
      if(_mystream_stream_oready) begin
        _tmp_565 <= _tmp_564;
      end 
      if(_tmp_551) begin
        _mystream_sum_vec8_sink_mode <= 5'b1;
        _mystream_sum_vec8_sink_offset <= _tmp_557;
        _mystream_sum_vec8_sink_size <= _tmp_565;
        _mystream_sum_vec8_sink_stride <= 1;
      end 
      if(_tmp_551) begin
        _mystream_sum_vec8_sink_sel <= 73;
      end 
      if(_mystream_sink_start && _mystream_sum_vec8_sink_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_sum_vec8_sink_offset_buf <= _mystream_sum_vec8_sink_offset;
        _mystream_sum_vec8_sink_size_buf <= _mystream_sum_vec8_sink_size;
        _mystream_sum_vec8_sink_stride_buf <= _mystream_sum_vec8_sink_stride;
      end 
      if((_mystream_sum_vec8_sink_fsm_72 == 1) && _mystream_stream_oready) begin
        _mystream_sum_vec8_sink_waddr <= _mystream_sum_vec8_sink_offset_buf - _mystream_sum_vec8_sink_stride_buf;
        _mystream_sum_vec8_sink_count <= _mystream_sum_vec8_sink_size_buf;
      end 
      if((_mystream_sum_vec8_sink_fsm_72 == 2) && _mystream_stream_oready) begin
        _mystream_sum_vec8_sink_waddr <= _mystream_sum_vec8_sink_waddr + _mystream_sum_vec8_sink_stride_buf;
        _mystream_sum_vec8_sink_wdata <= mystream_sum_vec8_data;
        _mystream_sum_vec8_sink_wenable <= 1;
        _mystream_sum_vec8_sink_count <= _mystream_sum_vec8_sink_count - 1;
      end 
      if(_mystream_stream_oready) begin
        _tmp_567 <= _set_flag_566;
      end 
      if(_mystream_stream_oready) begin
        _tmp_568 <= _tmp_567;
      end 
      if(_mystream_stream_oready) begin
        _tmp_569 <= _tmp_568;
      end 
      if(_mystream_stream_oready) begin
        _tmp_570 <= _tmp_569;
      end 
      if(_mystream_stream_oready) begin
        _tmp_571 <= _tmp_570;
      end 
      if(_mystream_stream_oready) begin
        _tmp_572 <= _tmp_571;
      end 
      if(_mystream_stream_oready) begin
        _tmp_573 <= _th_comp_offset_4;
      end 
      if(_mystream_stream_oready) begin
        _tmp_574 <= _tmp_573;
      end 
      if(_mystream_stream_oready) begin
        _tmp_575 <= _tmp_574;
      end 
      if(_mystream_stream_oready) begin
        _tmp_576 <= _tmp_575;
      end 
      if(_mystream_stream_oready) begin
        _tmp_577 <= _tmp_576;
      end 
      if(_mystream_stream_oready) begin
        _tmp_578 <= _tmp_577;
      end 
      if(_mystream_stream_oready) begin
        _tmp_581 <= _tmp_580;
      end 
      if(_mystream_stream_oready) begin
        _tmp_582 <= _tmp_581;
      end 
      if(_mystream_stream_oready) begin
        _tmp_583 <= _tmp_582;
      end 
      if(_mystream_stream_oready) begin
        _tmp_584 <= _tmp_583;
      end 
      if(_mystream_stream_oready) begin
        _tmp_585 <= _tmp_584;
      end 
      if(_mystream_stream_oready) begin
        _tmp_586 <= _tmp_585;
      end 
      if(_tmp_572) begin
        _mystream_sum_vec9_sink_mode <= 5'b1;
        _mystream_sum_vec9_sink_offset <= _tmp_578;
        _mystream_sum_vec9_sink_size <= _tmp_586;
        _mystream_sum_vec9_sink_stride <= 1;
      end 
      if(_tmp_572) begin
        _mystream_sum_vec9_sink_sel <= 74;
      end 
      if(_mystream_sink_start && _mystream_sum_vec9_sink_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_sum_vec9_sink_offset_buf <= _mystream_sum_vec9_sink_offset;
        _mystream_sum_vec9_sink_size_buf <= _mystream_sum_vec9_sink_size;
        _mystream_sum_vec9_sink_stride_buf <= _mystream_sum_vec9_sink_stride;
      end 
      if((_mystream_sum_vec9_sink_fsm_73 == 1) && _mystream_stream_oready) begin
        _mystream_sum_vec9_sink_waddr <= _mystream_sum_vec9_sink_offset_buf - _mystream_sum_vec9_sink_stride_buf;
        _mystream_sum_vec9_sink_count <= _mystream_sum_vec9_sink_size_buf;
      end 
      if((_mystream_sum_vec9_sink_fsm_73 == 2) && _mystream_stream_oready) begin
        _mystream_sum_vec9_sink_waddr <= _mystream_sum_vec9_sink_waddr + _mystream_sum_vec9_sink_stride_buf;
        _mystream_sum_vec9_sink_wdata <= mystream_sum_vec9_data;
        _mystream_sum_vec9_sink_wenable <= 1;
        _mystream_sum_vec9_sink_count <= _mystream_sum_vec9_sink_count - 1;
      end 
      if(_mystream_stream_oready) begin
        _tmp_588 <= _set_flag_587;
      end 
      if(_mystream_stream_oready) begin
        _tmp_589 <= _tmp_588;
      end 
      if(_mystream_stream_oready) begin
        _tmp_590 <= _tmp_589;
      end 
      if(_mystream_stream_oready) begin
        _tmp_591 <= _tmp_590;
      end 
      if(_mystream_stream_oready) begin
        _tmp_592 <= _tmp_591;
      end 
      if(_mystream_stream_oready) begin
        _tmp_593 <= _tmp_592;
      end 
      if(_mystream_stream_oready) begin
        _tmp_594 <= _th_comp_offset_4;
      end 
      if(_mystream_stream_oready) begin
        _tmp_595 <= _tmp_594;
      end 
      if(_mystream_stream_oready) begin
        _tmp_596 <= _tmp_595;
      end 
      if(_mystream_stream_oready) begin
        _tmp_597 <= _tmp_596;
      end 
      if(_mystream_stream_oready) begin
        _tmp_598 <= _tmp_597;
      end 
      if(_mystream_stream_oready) begin
        _tmp_599 <= _tmp_598;
      end 
      if(_mystream_stream_oready) begin
        _tmp_602 <= _tmp_601;
      end 
      if(_mystream_stream_oready) begin
        _tmp_603 <= _tmp_602;
      end 
      if(_mystream_stream_oready) begin
        _tmp_604 <= _tmp_603;
      end 
      if(_mystream_stream_oready) begin
        _tmp_605 <= _tmp_604;
      end 
      if(_mystream_stream_oready) begin
        _tmp_606 <= _tmp_605;
      end 
      if(_mystream_stream_oready) begin
        _tmp_607 <= _tmp_606;
      end 
      if(_tmp_593) begin
        _mystream_sum_vec10_sink_mode <= 5'b1;
        _mystream_sum_vec10_sink_offset <= _tmp_599;
        _mystream_sum_vec10_sink_size <= _tmp_607;
        _mystream_sum_vec10_sink_stride <= 1;
      end 
      if(_tmp_593) begin
        _mystream_sum_vec10_sink_sel <= 75;
      end 
      if(_mystream_sink_start && _mystream_sum_vec10_sink_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_sum_vec10_sink_offset_buf <= _mystream_sum_vec10_sink_offset;
        _mystream_sum_vec10_sink_size_buf <= _mystream_sum_vec10_sink_size;
        _mystream_sum_vec10_sink_stride_buf <= _mystream_sum_vec10_sink_stride;
      end 
      if((_mystream_sum_vec10_sink_fsm_74 == 1) && _mystream_stream_oready) begin
        _mystream_sum_vec10_sink_waddr <= _mystream_sum_vec10_sink_offset_buf - _mystream_sum_vec10_sink_stride_buf;
        _mystream_sum_vec10_sink_count <= _mystream_sum_vec10_sink_size_buf;
      end 
      if((_mystream_sum_vec10_sink_fsm_74 == 2) && _mystream_stream_oready) begin
        _mystream_sum_vec10_sink_waddr <= _mystream_sum_vec10_sink_waddr + _mystream_sum_vec10_sink_stride_buf;
        _mystream_sum_vec10_sink_wdata <= mystream_sum_vec10_data;
        _mystream_sum_vec10_sink_wenable <= 1;
        _mystream_sum_vec10_sink_count <= _mystream_sum_vec10_sink_count - 1;
      end 
      if(_mystream_stream_oready) begin
        _tmp_609 <= _set_flag_608;
      end 
      if(_mystream_stream_oready) begin
        _tmp_610 <= _tmp_609;
      end 
      if(_mystream_stream_oready) begin
        _tmp_611 <= _tmp_610;
      end 
      if(_mystream_stream_oready) begin
        _tmp_612 <= _tmp_611;
      end 
      if(_mystream_stream_oready) begin
        _tmp_613 <= _tmp_612;
      end 
      if(_mystream_stream_oready) begin
        _tmp_614 <= _tmp_613;
      end 
      if(_mystream_stream_oready) begin
        _tmp_615 <= _th_comp_offset_4;
      end 
      if(_mystream_stream_oready) begin
        _tmp_616 <= _tmp_615;
      end 
      if(_mystream_stream_oready) begin
        _tmp_617 <= _tmp_616;
      end 
      if(_mystream_stream_oready) begin
        _tmp_618 <= _tmp_617;
      end 
      if(_mystream_stream_oready) begin
        _tmp_619 <= _tmp_618;
      end 
      if(_mystream_stream_oready) begin
        _tmp_620 <= _tmp_619;
      end 
      if(_mystream_stream_oready) begin
        _tmp_623 <= _tmp_622;
      end 
      if(_mystream_stream_oready) begin
        _tmp_624 <= _tmp_623;
      end 
      if(_mystream_stream_oready) begin
        _tmp_625 <= _tmp_624;
      end 
      if(_mystream_stream_oready) begin
        _tmp_626 <= _tmp_625;
      end 
      if(_mystream_stream_oready) begin
        _tmp_627 <= _tmp_626;
      end 
      if(_mystream_stream_oready) begin
        _tmp_628 <= _tmp_627;
      end 
      if(_tmp_614) begin
        _mystream_sum_vec11_sink_mode <= 5'b1;
        _mystream_sum_vec11_sink_offset <= _tmp_620;
        _mystream_sum_vec11_sink_size <= _tmp_628;
        _mystream_sum_vec11_sink_stride <= 1;
      end 
      if(_tmp_614) begin
        _mystream_sum_vec11_sink_sel <= 76;
      end 
      if(_mystream_sink_start && _mystream_sum_vec11_sink_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_sum_vec11_sink_offset_buf <= _mystream_sum_vec11_sink_offset;
        _mystream_sum_vec11_sink_size_buf <= _mystream_sum_vec11_sink_size;
        _mystream_sum_vec11_sink_stride_buf <= _mystream_sum_vec11_sink_stride;
      end 
      if((_mystream_sum_vec11_sink_fsm_75 == 1) && _mystream_stream_oready) begin
        _mystream_sum_vec11_sink_waddr <= _mystream_sum_vec11_sink_offset_buf - _mystream_sum_vec11_sink_stride_buf;
        _mystream_sum_vec11_sink_count <= _mystream_sum_vec11_sink_size_buf;
      end 
      if((_mystream_sum_vec11_sink_fsm_75 == 2) && _mystream_stream_oready) begin
        _mystream_sum_vec11_sink_waddr <= _mystream_sum_vec11_sink_waddr + _mystream_sum_vec11_sink_stride_buf;
        _mystream_sum_vec11_sink_wdata <= mystream_sum_vec11_data;
        _mystream_sum_vec11_sink_wenable <= 1;
        _mystream_sum_vec11_sink_count <= _mystream_sum_vec11_sink_count - 1;
      end 
      if(_mystream_stream_oready) begin
        _tmp_630 <= _set_flag_629;
      end 
      if(_mystream_stream_oready) begin
        _tmp_631 <= _tmp_630;
      end 
      if(_mystream_stream_oready) begin
        _tmp_632 <= _tmp_631;
      end 
      if(_mystream_stream_oready) begin
        _tmp_633 <= _tmp_632;
      end 
      if(_mystream_stream_oready) begin
        _tmp_634 <= _tmp_633;
      end 
      if(_mystream_stream_oready) begin
        _tmp_635 <= _tmp_634;
      end 
      if(_mystream_stream_oready) begin
        _tmp_636 <= _th_comp_offset_4;
      end 
      if(_mystream_stream_oready) begin
        _tmp_637 <= _tmp_636;
      end 
      if(_mystream_stream_oready) begin
        _tmp_638 <= _tmp_637;
      end 
      if(_mystream_stream_oready) begin
        _tmp_639 <= _tmp_638;
      end 
      if(_mystream_stream_oready) begin
        _tmp_640 <= _tmp_639;
      end 
      if(_mystream_stream_oready) begin
        _tmp_641 <= _tmp_640;
      end 
      if(_mystream_stream_oready) begin
        _tmp_644 <= _tmp_643;
      end 
      if(_mystream_stream_oready) begin
        _tmp_645 <= _tmp_644;
      end 
      if(_mystream_stream_oready) begin
        _tmp_646 <= _tmp_645;
      end 
      if(_mystream_stream_oready) begin
        _tmp_647 <= _tmp_646;
      end 
      if(_mystream_stream_oready) begin
        _tmp_648 <= _tmp_647;
      end 
      if(_mystream_stream_oready) begin
        _tmp_649 <= _tmp_648;
      end 
      if(_tmp_635) begin
        _mystream_sum_vec12_sink_mode <= 5'b1;
        _mystream_sum_vec12_sink_offset <= _tmp_641;
        _mystream_sum_vec12_sink_size <= _tmp_649;
        _mystream_sum_vec12_sink_stride <= 1;
      end 
      if(_tmp_635) begin
        _mystream_sum_vec12_sink_sel <= 77;
      end 
      if(_mystream_sink_start && _mystream_sum_vec12_sink_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_sum_vec12_sink_offset_buf <= _mystream_sum_vec12_sink_offset;
        _mystream_sum_vec12_sink_size_buf <= _mystream_sum_vec12_sink_size;
        _mystream_sum_vec12_sink_stride_buf <= _mystream_sum_vec12_sink_stride;
      end 
      if((_mystream_sum_vec12_sink_fsm_76 == 1) && _mystream_stream_oready) begin
        _mystream_sum_vec12_sink_waddr <= _mystream_sum_vec12_sink_offset_buf - _mystream_sum_vec12_sink_stride_buf;
        _mystream_sum_vec12_sink_count <= _mystream_sum_vec12_sink_size_buf;
      end 
      if((_mystream_sum_vec12_sink_fsm_76 == 2) && _mystream_stream_oready) begin
        _mystream_sum_vec12_sink_waddr <= _mystream_sum_vec12_sink_waddr + _mystream_sum_vec12_sink_stride_buf;
        _mystream_sum_vec12_sink_wdata <= mystream_sum_vec12_data;
        _mystream_sum_vec12_sink_wenable <= 1;
        _mystream_sum_vec12_sink_count <= _mystream_sum_vec12_sink_count - 1;
      end 
      if(_mystream_stream_oready) begin
        _tmp_651 <= _set_flag_650;
      end 
      if(_mystream_stream_oready) begin
        _tmp_652 <= _tmp_651;
      end 
      if(_mystream_stream_oready) begin
        _tmp_653 <= _tmp_652;
      end 
      if(_mystream_stream_oready) begin
        _tmp_654 <= _tmp_653;
      end 
      if(_mystream_stream_oready) begin
        _tmp_655 <= _tmp_654;
      end 
      if(_mystream_stream_oready) begin
        _tmp_656 <= _tmp_655;
      end 
      if(_mystream_stream_oready) begin
        _tmp_657 <= _th_comp_offset_4;
      end 
      if(_mystream_stream_oready) begin
        _tmp_658 <= _tmp_657;
      end 
      if(_mystream_stream_oready) begin
        _tmp_659 <= _tmp_658;
      end 
      if(_mystream_stream_oready) begin
        _tmp_660 <= _tmp_659;
      end 
      if(_mystream_stream_oready) begin
        _tmp_661 <= _tmp_660;
      end 
      if(_mystream_stream_oready) begin
        _tmp_662 <= _tmp_661;
      end 
      if(_mystream_stream_oready) begin
        _tmp_665 <= _tmp_664;
      end 
      if(_mystream_stream_oready) begin
        _tmp_666 <= _tmp_665;
      end 
      if(_mystream_stream_oready) begin
        _tmp_667 <= _tmp_666;
      end 
      if(_mystream_stream_oready) begin
        _tmp_668 <= _tmp_667;
      end 
      if(_mystream_stream_oready) begin
        _tmp_669 <= _tmp_668;
      end 
      if(_mystream_stream_oready) begin
        _tmp_670 <= _tmp_669;
      end 
      if(_tmp_656) begin
        _mystream_sum_vec13_sink_mode <= 5'b1;
        _mystream_sum_vec13_sink_offset <= _tmp_662;
        _mystream_sum_vec13_sink_size <= _tmp_670;
        _mystream_sum_vec13_sink_stride <= 1;
      end 
      if(_tmp_656) begin
        _mystream_sum_vec13_sink_sel <= 78;
      end 
      if(_mystream_sink_start && _mystream_sum_vec13_sink_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_sum_vec13_sink_offset_buf <= _mystream_sum_vec13_sink_offset;
        _mystream_sum_vec13_sink_size_buf <= _mystream_sum_vec13_sink_size;
        _mystream_sum_vec13_sink_stride_buf <= _mystream_sum_vec13_sink_stride;
      end 
      if((_mystream_sum_vec13_sink_fsm_77 == 1) && _mystream_stream_oready) begin
        _mystream_sum_vec13_sink_waddr <= _mystream_sum_vec13_sink_offset_buf - _mystream_sum_vec13_sink_stride_buf;
        _mystream_sum_vec13_sink_count <= _mystream_sum_vec13_sink_size_buf;
      end 
      if((_mystream_sum_vec13_sink_fsm_77 == 2) && _mystream_stream_oready) begin
        _mystream_sum_vec13_sink_waddr <= _mystream_sum_vec13_sink_waddr + _mystream_sum_vec13_sink_stride_buf;
        _mystream_sum_vec13_sink_wdata <= mystream_sum_vec13_data;
        _mystream_sum_vec13_sink_wenable <= 1;
        _mystream_sum_vec13_sink_count <= _mystream_sum_vec13_sink_count - 1;
      end 
      if(_mystream_stream_oready) begin
        _tmp_672 <= _set_flag_671;
      end 
      if(_mystream_stream_oready) begin
        _tmp_673 <= _tmp_672;
      end 
      if(_mystream_stream_oready) begin
        _tmp_674 <= _tmp_673;
      end 
      if(_mystream_stream_oready) begin
        _tmp_675 <= _tmp_674;
      end 
      if(_mystream_stream_oready) begin
        _tmp_676 <= _tmp_675;
      end 
      if(_mystream_stream_oready) begin
        _tmp_677 <= _tmp_676;
      end 
      if(_mystream_stream_oready) begin
        _tmp_678 <= _th_comp_offset_4;
      end 
      if(_mystream_stream_oready) begin
        _tmp_679 <= _tmp_678;
      end 
      if(_mystream_stream_oready) begin
        _tmp_680 <= _tmp_679;
      end 
      if(_mystream_stream_oready) begin
        _tmp_681 <= _tmp_680;
      end 
      if(_mystream_stream_oready) begin
        _tmp_682 <= _tmp_681;
      end 
      if(_mystream_stream_oready) begin
        _tmp_683 <= _tmp_682;
      end 
      if(_mystream_stream_oready) begin
        _tmp_686 <= _tmp_685;
      end 
      if(_mystream_stream_oready) begin
        _tmp_687 <= _tmp_686;
      end 
      if(_mystream_stream_oready) begin
        _tmp_688 <= _tmp_687;
      end 
      if(_mystream_stream_oready) begin
        _tmp_689 <= _tmp_688;
      end 
      if(_mystream_stream_oready) begin
        _tmp_690 <= _tmp_689;
      end 
      if(_mystream_stream_oready) begin
        _tmp_691 <= _tmp_690;
      end 
      if(_tmp_677) begin
        _mystream_sum_vec14_sink_mode <= 5'b1;
        _mystream_sum_vec14_sink_offset <= _tmp_683;
        _mystream_sum_vec14_sink_size <= _tmp_691;
        _mystream_sum_vec14_sink_stride <= 1;
      end 
      if(_tmp_677) begin
        _mystream_sum_vec14_sink_sel <= 79;
      end 
      if(_mystream_sink_start && _mystream_sum_vec14_sink_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_sum_vec14_sink_offset_buf <= _mystream_sum_vec14_sink_offset;
        _mystream_sum_vec14_sink_size_buf <= _mystream_sum_vec14_sink_size;
        _mystream_sum_vec14_sink_stride_buf <= _mystream_sum_vec14_sink_stride;
      end 
      if((_mystream_sum_vec14_sink_fsm_78 == 1) && _mystream_stream_oready) begin
        _mystream_sum_vec14_sink_waddr <= _mystream_sum_vec14_sink_offset_buf - _mystream_sum_vec14_sink_stride_buf;
        _mystream_sum_vec14_sink_count <= _mystream_sum_vec14_sink_size_buf;
      end 
      if((_mystream_sum_vec14_sink_fsm_78 == 2) && _mystream_stream_oready) begin
        _mystream_sum_vec14_sink_waddr <= _mystream_sum_vec14_sink_waddr + _mystream_sum_vec14_sink_stride_buf;
        _mystream_sum_vec14_sink_wdata <= mystream_sum_vec14_data;
        _mystream_sum_vec14_sink_wenable <= 1;
        _mystream_sum_vec14_sink_count <= _mystream_sum_vec14_sink_count - 1;
      end 
      if(_mystream_stream_oready) begin
        _tmp_693 <= _set_flag_692;
      end 
      if(_mystream_stream_oready) begin
        _tmp_694 <= _tmp_693;
      end 
      if(_mystream_stream_oready) begin
        _tmp_695 <= _tmp_694;
      end 
      if(_mystream_stream_oready) begin
        _tmp_696 <= _tmp_695;
      end 
      if(_mystream_stream_oready) begin
        _tmp_697 <= _tmp_696;
      end 
      if(_mystream_stream_oready) begin
        _tmp_698 <= _tmp_697;
      end 
      if(_mystream_stream_oready) begin
        _tmp_699 <= _th_comp_offset_4;
      end 
      if(_mystream_stream_oready) begin
        _tmp_700 <= _tmp_699;
      end 
      if(_mystream_stream_oready) begin
        _tmp_701 <= _tmp_700;
      end 
      if(_mystream_stream_oready) begin
        _tmp_702 <= _tmp_701;
      end 
      if(_mystream_stream_oready) begin
        _tmp_703 <= _tmp_702;
      end 
      if(_mystream_stream_oready) begin
        _tmp_704 <= _tmp_703;
      end 
      if(_mystream_stream_oready) begin
        _tmp_707 <= _tmp_706;
      end 
      if(_mystream_stream_oready) begin
        _tmp_708 <= _tmp_707;
      end 
      if(_mystream_stream_oready) begin
        _tmp_709 <= _tmp_708;
      end 
      if(_mystream_stream_oready) begin
        _tmp_710 <= _tmp_709;
      end 
      if(_mystream_stream_oready) begin
        _tmp_711 <= _tmp_710;
      end 
      if(_mystream_stream_oready) begin
        _tmp_712 <= _tmp_711;
      end 
      if(_tmp_698) begin
        _mystream_sum_vec15_sink_mode <= 5'b1;
        _mystream_sum_vec15_sink_offset <= _tmp_704;
        _mystream_sum_vec15_sink_size <= _tmp_712;
        _mystream_sum_vec15_sink_stride <= 1;
      end 
      if(_tmp_698) begin
        _mystream_sum_vec15_sink_sel <= 80;
      end 
      if(_mystream_sink_start && _mystream_sum_vec15_sink_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_sum_vec15_sink_offset_buf <= _mystream_sum_vec15_sink_offset;
        _mystream_sum_vec15_sink_size_buf <= _mystream_sum_vec15_sink_size;
        _mystream_sum_vec15_sink_stride_buf <= _mystream_sum_vec15_sink_stride;
      end 
      if((_mystream_sum_vec15_sink_fsm_79 == 1) && _mystream_stream_oready) begin
        _mystream_sum_vec15_sink_waddr <= _mystream_sum_vec15_sink_offset_buf - _mystream_sum_vec15_sink_stride_buf;
        _mystream_sum_vec15_sink_count <= _mystream_sum_vec15_sink_size_buf;
      end 
      if((_mystream_sum_vec15_sink_fsm_79 == 2) && _mystream_stream_oready) begin
        _mystream_sum_vec15_sink_waddr <= _mystream_sum_vec15_sink_waddr + _mystream_sum_vec15_sink_stride_buf;
        _mystream_sum_vec15_sink_wdata <= mystream_sum_vec15_data;
        _mystream_sum_vec15_sink_wenable <= 1;
        _mystream_sum_vec15_sink_count <= _mystream_sum_vec15_sink_count - 1;
      end 
      if(_mystream_stream_oready) begin
        _tmp_714 <= _set_flag_713;
      end 
      if(_mystream_stream_oready) begin
        _tmp_715 <= _tmp_714;
      end 
      if(_mystream_stream_oready) begin
        _tmp_716 <= _tmp_715;
      end 
      if(_mystream_stream_oready) begin
        _tmp_717 <= _tmp_716;
      end 
      if(_mystream_stream_oready) begin
        _tmp_718 <= _tmp_717;
      end 
      if(_mystream_stream_oready) begin
        _tmp_719 <= _tmp_718;
      end 
      if(_mystream_stream_oready) begin
        _tmp_720 <= _th_comp_offset_4;
      end 
      if(_mystream_stream_oready) begin
        _tmp_721 <= _tmp_720;
      end 
      if(_mystream_stream_oready) begin
        _tmp_722 <= _tmp_721;
      end 
      if(_mystream_stream_oready) begin
        _tmp_723 <= _tmp_722;
      end 
      if(_mystream_stream_oready) begin
        _tmp_724 <= _tmp_723;
      end 
      if(_mystream_stream_oready) begin
        _tmp_725 <= _tmp_724;
      end 
      if(_mystream_stream_oready) begin
        _tmp_728 <= _tmp_727;
      end 
      if(_mystream_stream_oready) begin
        _tmp_729 <= _tmp_728;
      end 
      if(_mystream_stream_oready) begin
        _tmp_730 <= _tmp_729;
      end 
      if(_mystream_stream_oready) begin
        _tmp_731 <= _tmp_730;
      end 
      if(_mystream_stream_oready) begin
        _tmp_732 <= _tmp_731;
      end 
      if(_mystream_stream_oready) begin
        _tmp_733 <= _tmp_732;
      end 
      if(_tmp_719) begin
        _mystream_sum_vec16_sink_mode <= 5'b1;
        _mystream_sum_vec16_sink_offset <= _tmp_725;
        _mystream_sum_vec16_sink_size <= _tmp_733;
        _mystream_sum_vec16_sink_stride <= 1;
      end 
      if(_tmp_719) begin
        _mystream_sum_vec16_sink_sel <= 81;
      end 
      if(_mystream_sink_start && _mystream_sum_vec16_sink_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_sum_vec16_sink_offset_buf <= _mystream_sum_vec16_sink_offset;
        _mystream_sum_vec16_sink_size_buf <= _mystream_sum_vec16_sink_size;
        _mystream_sum_vec16_sink_stride_buf <= _mystream_sum_vec16_sink_stride;
      end 
      if((_mystream_sum_vec16_sink_fsm_80 == 1) && _mystream_stream_oready) begin
        _mystream_sum_vec16_sink_waddr <= _mystream_sum_vec16_sink_offset_buf - _mystream_sum_vec16_sink_stride_buf;
        _mystream_sum_vec16_sink_count <= _mystream_sum_vec16_sink_size_buf;
      end 
      if((_mystream_sum_vec16_sink_fsm_80 == 2) && _mystream_stream_oready) begin
        _mystream_sum_vec16_sink_waddr <= _mystream_sum_vec16_sink_waddr + _mystream_sum_vec16_sink_stride_buf;
        _mystream_sum_vec16_sink_wdata <= mystream_sum_vec16_data;
        _mystream_sum_vec16_sink_wenable <= 1;
        _mystream_sum_vec16_sink_count <= _mystream_sum_vec16_sink_count - 1;
      end 
      if(_mystream_stream_oready) begin
        _tmp_735 <= _set_flag_734;
      end 
      if(_mystream_stream_oready) begin
        _tmp_736 <= _tmp_735;
      end 
      if(_mystream_stream_oready) begin
        _tmp_737 <= _tmp_736;
      end 
      if(_mystream_stream_oready) begin
        _tmp_738 <= _tmp_737;
      end 
      if(_mystream_stream_oready) begin
        _tmp_739 <= _tmp_738;
      end 
      if(_mystream_stream_oready) begin
        _tmp_740 <= _tmp_739;
      end 
      if(_mystream_stream_oready) begin
        _tmp_741 <= _th_comp_offset_4;
      end 
      if(_mystream_stream_oready) begin
        _tmp_742 <= _tmp_741;
      end 
      if(_mystream_stream_oready) begin
        _tmp_743 <= _tmp_742;
      end 
      if(_mystream_stream_oready) begin
        _tmp_744 <= _tmp_743;
      end 
      if(_mystream_stream_oready) begin
        _tmp_745 <= _tmp_744;
      end 
      if(_mystream_stream_oready) begin
        _tmp_746 <= _tmp_745;
      end 
      if(_mystream_stream_oready) begin
        _tmp_749 <= _tmp_748;
      end 
      if(_mystream_stream_oready) begin
        _tmp_750 <= _tmp_749;
      end 
      if(_mystream_stream_oready) begin
        _tmp_751 <= _tmp_750;
      end 
      if(_mystream_stream_oready) begin
        _tmp_752 <= _tmp_751;
      end 
      if(_mystream_stream_oready) begin
        _tmp_753 <= _tmp_752;
      end 
      if(_mystream_stream_oready) begin
        _tmp_754 <= _tmp_753;
      end 
      if(_tmp_740) begin
        _mystream_sum_vec17_sink_mode <= 5'b1;
        _mystream_sum_vec17_sink_offset <= _tmp_746;
        _mystream_sum_vec17_sink_size <= _tmp_754;
        _mystream_sum_vec17_sink_stride <= 1;
      end 
      if(_tmp_740) begin
        _mystream_sum_vec17_sink_sel <= 82;
      end 
      if(_mystream_sink_start && _mystream_sum_vec17_sink_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_sum_vec17_sink_offset_buf <= _mystream_sum_vec17_sink_offset;
        _mystream_sum_vec17_sink_size_buf <= _mystream_sum_vec17_sink_size;
        _mystream_sum_vec17_sink_stride_buf <= _mystream_sum_vec17_sink_stride;
      end 
      if((_mystream_sum_vec17_sink_fsm_81 == 1) && _mystream_stream_oready) begin
        _mystream_sum_vec17_sink_waddr <= _mystream_sum_vec17_sink_offset_buf - _mystream_sum_vec17_sink_stride_buf;
        _mystream_sum_vec17_sink_count <= _mystream_sum_vec17_sink_size_buf;
      end 
      if((_mystream_sum_vec17_sink_fsm_81 == 2) && _mystream_stream_oready) begin
        _mystream_sum_vec17_sink_waddr <= _mystream_sum_vec17_sink_waddr + _mystream_sum_vec17_sink_stride_buf;
        _mystream_sum_vec17_sink_wdata <= mystream_sum_vec17_data;
        _mystream_sum_vec17_sink_wenable <= 1;
        _mystream_sum_vec17_sink_count <= _mystream_sum_vec17_sink_count - 1;
      end 
      if(_mystream_stream_oready) begin
        _tmp_756 <= _set_flag_755;
      end 
      if(_mystream_stream_oready) begin
        _tmp_757 <= _tmp_756;
      end 
      if(_mystream_stream_oready) begin
        _tmp_758 <= _tmp_757;
      end 
      if(_mystream_stream_oready) begin
        _tmp_759 <= _tmp_758;
      end 
      if(_mystream_stream_oready) begin
        _tmp_760 <= _tmp_759;
      end 
      if(_mystream_stream_oready) begin
        _tmp_761 <= _tmp_760;
      end 
      if(_mystream_stream_oready) begin
        _tmp_762 <= _th_comp_offset_4;
      end 
      if(_mystream_stream_oready) begin
        _tmp_763 <= _tmp_762;
      end 
      if(_mystream_stream_oready) begin
        _tmp_764 <= _tmp_763;
      end 
      if(_mystream_stream_oready) begin
        _tmp_765 <= _tmp_764;
      end 
      if(_mystream_stream_oready) begin
        _tmp_766 <= _tmp_765;
      end 
      if(_mystream_stream_oready) begin
        _tmp_767 <= _tmp_766;
      end 
      if(_mystream_stream_oready) begin
        _tmp_770 <= _tmp_769;
      end 
      if(_mystream_stream_oready) begin
        _tmp_771 <= _tmp_770;
      end 
      if(_mystream_stream_oready) begin
        _tmp_772 <= _tmp_771;
      end 
      if(_mystream_stream_oready) begin
        _tmp_773 <= _tmp_772;
      end 
      if(_mystream_stream_oready) begin
        _tmp_774 <= _tmp_773;
      end 
      if(_mystream_stream_oready) begin
        _tmp_775 <= _tmp_774;
      end 
      if(_tmp_761) begin
        _mystream_sum_vec18_sink_mode <= 5'b1;
        _mystream_sum_vec18_sink_offset <= _tmp_767;
        _mystream_sum_vec18_sink_size <= _tmp_775;
        _mystream_sum_vec18_sink_stride <= 1;
      end 
      if(_tmp_761) begin
        _mystream_sum_vec18_sink_sel <= 83;
      end 
      if(_mystream_sink_start && _mystream_sum_vec18_sink_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_sum_vec18_sink_offset_buf <= _mystream_sum_vec18_sink_offset;
        _mystream_sum_vec18_sink_size_buf <= _mystream_sum_vec18_sink_size;
        _mystream_sum_vec18_sink_stride_buf <= _mystream_sum_vec18_sink_stride;
      end 
      if((_mystream_sum_vec18_sink_fsm_82 == 1) && _mystream_stream_oready) begin
        _mystream_sum_vec18_sink_waddr <= _mystream_sum_vec18_sink_offset_buf - _mystream_sum_vec18_sink_stride_buf;
        _mystream_sum_vec18_sink_count <= _mystream_sum_vec18_sink_size_buf;
      end 
      if((_mystream_sum_vec18_sink_fsm_82 == 2) && _mystream_stream_oready) begin
        _mystream_sum_vec18_sink_waddr <= _mystream_sum_vec18_sink_waddr + _mystream_sum_vec18_sink_stride_buf;
        _mystream_sum_vec18_sink_wdata <= mystream_sum_vec18_data;
        _mystream_sum_vec18_sink_wenable <= 1;
        _mystream_sum_vec18_sink_count <= _mystream_sum_vec18_sink_count - 1;
      end 
      if(_mystream_stream_oready) begin
        _tmp_777 <= _set_flag_776;
      end 
      if(_mystream_stream_oready) begin
        _tmp_778 <= _tmp_777;
      end 
      if(_mystream_stream_oready) begin
        _tmp_779 <= _tmp_778;
      end 
      if(_mystream_stream_oready) begin
        _tmp_780 <= _tmp_779;
      end 
      if(_mystream_stream_oready) begin
        _tmp_781 <= _tmp_780;
      end 
      if(_mystream_stream_oready) begin
        _tmp_782 <= _tmp_781;
      end 
      if(_mystream_stream_oready) begin
        _tmp_783 <= _th_comp_offset_4;
      end 
      if(_mystream_stream_oready) begin
        _tmp_784 <= _tmp_783;
      end 
      if(_mystream_stream_oready) begin
        _tmp_785 <= _tmp_784;
      end 
      if(_mystream_stream_oready) begin
        _tmp_786 <= _tmp_785;
      end 
      if(_mystream_stream_oready) begin
        _tmp_787 <= _tmp_786;
      end 
      if(_mystream_stream_oready) begin
        _tmp_788 <= _tmp_787;
      end 
      if(_mystream_stream_oready) begin
        _tmp_791 <= _tmp_790;
      end 
      if(_mystream_stream_oready) begin
        _tmp_792 <= _tmp_791;
      end 
      if(_mystream_stream_oready) begin
        _tmp_793 <= _tmp_792;
      end 
      if(_mystream_stream_oready) begin
        _tmp_794 <= _tmp_793;
      end 
      if(_mystream_stream_oready) begin
        _tmp_795 <= _tmp_794;
      end 
      if(_mystream_stream_oready) begin
        _tmp_796 <= _tmp_795;
      end 
      if(_tmp_782) begin
        _mystream_sum_vec19_sink_mode <= 5'b1;
        _mystream_sum_vec19_sink_offset <= _tmp_788;
        _mystream_sum_vec19_sink_size <= _tmp_796;
        _mystream_sum_vec19_sink_stride <= 1;
      end 
      if(_tmp_782) begin
        _mystream_sum_vec19_sink_sel <= 84;
      end 
      if(_mystream_sink_start && _mystream_sum_vec19_sink_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_sum_vec19_sink_offset_buf <= _mystream_sum_vec19_sink_offset;
        _mystream_sum_vec19_sink_size_buf <= _mystream_sum_vec19_sink_size;
        _mystream_sum_vec19_sink_stride_buf <= _mystream_sum_vec19_sink_stride;
      end 
      if((_mystream_sum_vec19_sink_fsm_83 == 1) && _mystream_stream_oready) begin
        _mystream_sum_vec19_sink_waddr <= _mystream_sum_vec19_sink_offset_buf - _mystream_sum_vec19_sink_stride_buf;
        _mystream_sum_vec19_sink_count <= _mystream_sum_vec19_sink_size_buf;
      end 
      if((_mystream_sum_vec19_sink_fsm_83 == 2) && _mystream_stream_oready) begin
        _mystream_sum_vec19_sink_waddr <= _mystream_sum_vec19_sink_waddr + _mystream_sum_vec19_sink_stride_buf;
        _mystream_sum_vec19_sink_wdata <= mystream_sum_vec19_data;
        _mystream_sum_vec19_sink_wenable <= 1;
        _mystream_sum_vec19_sink_count <= _mystream_sum_vec19_sink_count - 1;
      end 
      if(_mystream_stream_oready) begin
        _tmp_798 <= _set_flag_797;
      end 
      if(_mystream_stream_oready) begin
        _tmp_799 <= _tmp_798;
      end 
      if(_mystream_stream_oready) begin
        _tmp_800 <= _tmp_799;
      end 
      if(_mystream_stream_oready) begin
        _tmp_801 <= _tmp_800;
      end 
      if(_mystream_stream_oready) begin
        _tmp_802 <= _tmp_801;
      end 
      if(_mystream_stream_oready) begin
        _tmp_803 <= _tmp_802;
      end 
      if(_mystream_stream_oready) begin
        _tmp_804 <= _th_comp_offset_4;
      end 
      if(_mystream_stream_oready) begin
        _tmp_805 <= _tmp_804;
      end 
      if(_mystream_stream_oready) begin
        _tmp_806 <= _tmp_805;
      end 
      if(_mystream_stream_oready) begin
        _tmp_807 <= _tmp_806;
      end 
      if(_mystream_stream_oready) begin
        _tmp_808 <= _tmp_807;
      end 
      if(_mystream_stream_oready) begin
        _tmp_809 <= _tmp_808;
      end 
      if(_mystream_stream_oready) begin
        _tmp_812 <= _tmp_811;
      end 
      if(_mystream_stream_oready) begin
        _tmp_813 <= _tmp_812;
      end 
      if(_mystream_stream_oready) begin
        _tmp_814 <= _tmp_813;
      end 
      if(_mystream_stream_oready) begin
        _tmp_815 <= _tmp_814;
      end 
      if(_mystream_stream_oready) begin
        _tmp_816 <= _tmp_815;
      end 
      if(_mystream_stream_oready) begin
        _tmp_817 <= _tmp_816;
      end 
      if(_tmp_803) begin
        _mystream_sum_vec20_sink_mode <= 5'b1;
        _mystream_sum_vec20_sink_offset <= _tmp_809;
        _mystream_sum_vec20_sink_size <= _tmp_817;
        _mystream_sum_vec20_sink_stride <= 1;
      end 
      if(_tmp_803) begin
        _mystream_sum_vec20_sink_sel <= 85;
      end 
      if(_mystream_sink_start && _mystream_sum_vec20_sink_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_sum_vec20_sink_offset_buf <= _mystream_sum_vec20_sink_offset;
        _mystream_sum_vec20_sink_size_buf <= _mystream_sum_vec20_sink_size;
        _mystream_sum_vec20_sink_stride_buf <= _mystream_sum_vec20_sink_stride;
      end 
      if((_mystream_sum_vec20_sink_fsm_84 == 1) && _mystream_stream_oready) begin
        _mystream_sum_vec20_sink_waddr <= _mystream_sum_vec20_sink_offset_buf - _mystream_sum_vec20_sink_stride_buf;
        _mystream_sum_vec20_sink_count <= _mystream_sum_vec20_sink_size_buf;
      end 
      if((_mystream_sum_vec20_sink_fsm_84 == 2) && _mystream_stream_oready) begin
        _mystream_sum_vec20_sink_waddr <= _mystream_sum_vec20_sink_waddr + _mystream_sum_vec20_sink_stride_buf;
        _mystream_sum_vec20_sink_wdata <= mystream_sum_vec20_data;
        _mystream_sum_vec20_sink_wenable <= 1;
        _mystream_sum_vec20_sink_count <= _mystream_sum_vec20_sink_count - 1;
      end 
      if(_mystream_stream_oready) begin
        _tmp_819 <= _set_flag_818;
      end 
      if(_mystream_stream_oready) begin
        _tmp_820 <= _tmp_819;
      end 
      if(_mystream_stream_oready) begin
        _tmp_821 <= _tmp_820;
      end 
      if(_mystream_stream_oready) begin
        _tmp_822 <= _tmp_821;
      end 
      if(_mystream_stream_oready) begin
        _tmp_823 <= _tmp_822;
      end 
      if(_mystream_stream_oready) begin
        _tmp_824 <= _tmp_823;
      end 
      if(_mystream_stream_oready) begin
        _tmp_825 <= _th_comp_offset_4;
      end 
      if(_mystream_stream_oready) begin
        _tmp_826 <= _tmp_825;
      end 
      if(_mystream_stream_oready) begin
        _tmp_827 <= _tmp_826;
      end 
      if(_mystream_stream_oready) begin
        _tmp_828 <= _tmp_827;
      end 
      if(_mystream_stream_oready) begin
        _tmp_829 <= _tmp_828;
      end 
      if(_mystream_stream_oready) begin
        _tmp_830 <= _tmp_829;
      end 
      if(_mystream_stream_oready) begin
        _tmp_833 <= _tmp_832;
      end 
      if(_mystream_stream_oready) begin
        _tmp_834 <= _tmp_833;
      end 
      if(_mystream_stream_oready) begin
        _tmp_835 <= _tmp_834;
      end 
      if(_mystream_stream_oready) begin
        _tmp_836 <= _tmp_835;
      end 
      if(_mystream_stream_oready) begin
        _tmp_837 <= _tmp_836;
      end 
      if(_mystream_stream_oready) begin
        _tmp_838 <= _tmp_837;
      end 
      if(_tmp_824) begin
        _mystream_sum_vec21_sink_mode <= 5'b1;
        _mystream_sum_vec21_sink_offset <= _tmp_830;
        _mystream_sum_vec21_sink_size <= _tmp_838;
        _mystream_sum_vec21_sink_stride <= 1;
      end 
      if(_tmp_824) begin
        _mystream_sum_vec21_sink_sel <= 86;
      end 
      if(_mystream_sink_start && _mystream_sum_vec21_sink_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_sum_vec21_sink_offset_buf <= _mystream_sum_vec21_sink_offset;
        _mystream_sum_vec21_sink_size_buf <= _mystream_sum_vec21_sink_size;
        _mystream_sum_vec21_sink_stride_buf <= _mystream_sum_vec21_sink_stride;
      end 
      if((_mystream_sum_vec21_sink_fsm_85 == 1) && _mystream_stream_oready) begin
        _mystream_sum_vec21_sink_waddr <= _mystream_sum_vec21_sink_offset_buf - _mystream_sum_vec21_sink_stride_buf;
        _mystream_sum_vec21_sink_count <= _mystream_sum_vec21_sink_size_buf;
      end 
      if((_mystream_sum_vec21_sink_fsm_85 == 2) && _mystream_stream_oready) begin
        _mystream_sum_vec21_sink_waddr <= _mystream_sum_vec21_sink_waddr + _mystream_sum_vec21_sink_stride_buf;
        _mystream_sum_vec21_sink_wdata <= mystream_sum_vec21_data;
        _mystream_sum_vec21_sink_wenable <= 1;
        _mystream_sum_vec21_sink_count <= _mystream_sum_vec21_sink_count - 1;
      end 
      if(_mystream_stream_oready) begin
        _tmp_840 <= _set_flag_839;
      end 
      if(_mystream_stream_oready) begin
        _tmp_841 <= _tmp_840;
      end 
      if(_mystream_stream_oready) begin
        _tmp_842 <= _tmp_841;
      end 
      if(_mystream_stream_oready) begin
        _tmp_843 <= _tmp_842;
      end 
      if(_mystream_stream_oready) begin
        _tmp_844 <= _tmp_843;
      end 
      if(_mystream_stream_oready) begin
        _tmp_845 <= _tmp_844;
      end 
      if(_mystream_stream_oready) begin
        _tmp_846 <= _th_comp_offset_4;
      end 
      if(_mystream_stream_oready) begin
        _tmp_847 <= _tmp_846;
      end 
      if(_mystream_stream_oready) begin
        _tmp_848 <= _tmp_847;
      end 
      if(_mystream_stream_oready) begin
        _tmp_849 <= _tmp_848;
      end 
      if(_mystream_stream_oready) begin
        _tmp_850 <= _tmp_849;
      end 
      if(_mystream_stream_oready) begin
        _tmp_851 <= _tmp_850;
      end 
      if(_mystream_stream_oready) begin
        _tmp_854 <= _tmp_853;
      end 
      if(_mystream_stream_oready) begin
        _tmp_855 <= _tmp_854;
      end 
      if(_mystream_stream_oready) begin
        _tmp_856 <= _tmp_855;
      end 
      if(_mystream_stream_oready) begin
        _tmp_857 <= _tmp_856;
      end 
      if(_mystream_stream_oready) begin
        _tmp_858 <= _tmp_857;
      end 
      if(_mystream_stream_oready) begin
        _tmp_859 <= _tmp_858;
      end 
      if(_tmp_845) begin
        _mystream_sum_vec22_sink_mode <= 5'b1;
        _mystream_sum_vec22_sink_offset <= _tmp_851;
        _mystream_sum_vec22_sink_size <= _tmp_859;
        _mystream_sum_vec22_sink_stride <= 1;
      end 
      if(_tmp_845) begin
        _mystream_sum_vec22_sink_sel <= 87;
      end 
      if(_mystream_sink_start && _mystream_sum_vec22_sink_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_sum_vec22_sink_offset_buf <= _mystream_sum_vec22_sink_offset;
        _mystream_sum_vec22_sink_size_buf <= _mystream_sum_vec22_sink_size;
        _mystream_sum_vec22_sink_stride_buf <= _mystream_sum_vec22_sink_stride;
      end 
      if((_mystream_sum_vec22_sink_fsm_86 == 1) && _mystream_stream_oready) begin
        _mystream_sum_vec22_sink_waddr <= _mystream_sum_vec22_sink_offset_buf - _mystream_sum_vec22_sink_stride_buf;
        _mystream_sum_vec22_sink_count <= _mystream_sum_vec22_sink_size_buf;
      end 
      if((_mystream_sum_vec22_sink_fsm_86 == 2) && _mystream_stream_oready) begin
        _mystream_sum_vec22_sink_waddr <= _mystream_sum_vec22_sink_waddr + _mystream_sum_vec22_sink_stride_buf;
        _mystream_sum_vec22_sink_wdata <= mystream_sum_vec22_data;
        _mystream_sum_vec22_sink_wenable <= 1;
        _mystream_sum_vec22_sink_count <= _mystream_sum_vec22_sink_count - 1;
      end 
      if(_mystream_stream_oready) begin
        _tmp_861 <= _set_flag_860;
      end 
      if(_mystream_stream_oready) begin
        _tmp_862 <= _tmp_861;
      end 
      if(_mystream_stream_oready) begin
        _tmp_863 <= _tmp_862;
      end 
      if(_mystream_stream_oready) begin
        _tmp_864 <= _tmp_863;
      end 
      if(_mystream_stream_oready) begin
        _tmp_865 <= _tmp_864;
      end 
      if(_mystream_stream_oready) begin
        _tmp_866 <= _tmp_865;
      end 
      if(_mystream_stream_oready) begin
        _tmp_867 <= _th_comp_offset_4;
      end 
      if(_mystream_stream_oready) begin
        _tmp_868 <= _tmp_867;
      end 
      if(_mystream_stream_oready) begin
        _tmp_869 <= _tmp_868;
      end 
      if(_mystream_stream_oready) begin
        _tmp_870 <= _tmp_869;
      end 
      if(_mystream_stream_oready) begin
        _tmp_871 <= _tmp_870;
      end 
      if(_mystream_stream_oready) begin
        _tmp_872 <= _tmp_871;
      end 
      if(_mystream_stream_oready) begin
        _tmp_875 <= _tmp_874;
      end 
      if(_mystream_stream_oready) begin
        _tmp_876 <= _tmp_875;
      end 
      if(_mystream_stream_oready) begin
        _tmp_877 <= _tmp_876;
      end 
      if(_mystream_stream_oready) begin
        _tmp_878 <= _tmp_877;
      end 
      if(_mystream_stream_oready) begin
        _tmp_879 <= _tmp_878;
      end 
      if(_mystream_stream_oready) begin
        _tmp_880 <= _tmp_879;
      end 
      if(_tmp_866) begin
        _mystream_sum_vec23_sink_mode <= 5'b1;
        _mystream_sum_vec23_sink_offset <= _tmp_872;
        _mystream_sum_vec23_sink_size <= _tmp_880;
        _mystream_sum_vec23_sink_stride <= 1;
      end 
      if(_tmp_866) begin
        _mystream_sum_vec23_sink_sel <= 88;
      end 
      if(_mystream_sink_start && _mystream_sum_vec23_sink_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_sum_vec23_sink_offset_buf <= _mystream_sum_vec23_sink_offset;
        _mystream_sum_vec23_sink_size_buf <= _mystream_sum_vec23_sink_size;
        _mystream_sum_vec23_sink_stride_buf <= _mystream_sum_vec23_sink_stride;
      end 
      if((_mystream_sum_vec23_sink_fsm_87 == 1) && _mystream_stream_oready) begin
        _mystream_sum_vec23_sink_waddr <= _mystream_sum_vec23_sink_offset_buf - _mystream_sum_vec23_sink_stride_buf;
        _mystream_sum_vec23_sink_count <= _mystream_sum_vec23_sink_size_buf;
      end 
      if((_mystream_sum_vec23_sink_fsm_87 == 2) && _mystream_stream_oready) begin
        _mystream_sum_vec23_sink_waddr <= _mystream_sum_vec23_sink_waddr + _mystream_sum_vec23_sink_stride_buf;
        _mystream_sum_vec23_sink_wdata <= mystream_sum_vec23_data;
        _mystream_sum_vec23_sink_wenable <= 1;
        _mystream_sum_vec23_sink_count <= _mystream_sum_vec23_sink_count - 1;
      end 
      if(_mystream_stream_oready) begin
        _tmp_882 <= _set_flag_881;
      end 
      if(_mystream_stream_oready) begin
        _tmp_883 <= _tmp_882;
      end 
      if(_mystream_stream_oready) begin
        _tmp_884 <= _tmp_883;
      end 
      if(_mystream_stream_oready) begin
        _tmp_885 <= _tmp_884;
      end 
      if(_mystream_stream_oready) begin
        _tmp_886 <= _tmp_885;
      end 
      if(_mystream_stream_oready) begin
        _tmp_887 <= _tmp_886;
      end 
      if(_mystream_stream_oready) begin
        _tmp_888 <= _th_comp_offset_4;
      end 
      if(_mystream_stream_oready) begin
        _tmp_889 <= _tmp_888;
      end 
      if(_mystream_stream_oready) begin
        _tmp_890 <= _tmp_889;
      end 
      if(_mystream_stream_oready) begin
        _tmp_891 <= _tmp_890;
      end 
      if(_mystream_stream_oready) begin
        _tmp_892 <= _tmp_891;
      end 
      if(_mystream_stream_oready) begin
        _tmp_893 <= _tmp_892;
      end 
      if(_mystream_stream_oready) begin
        _tmp_896 <= _tmp_895;
      end 
      if(_mystream_stream_oready) begin
        _tmp_897 <= _tmp_896;
      end 
      if(_mystream_stream_oready) begin
        _tmp_898 <= _tmp_897;
      end 
      if(_mystream_stream_oready) begin
        _tmp_899 <= _tmp_898;
      end 
      if(_mystream_stream_oready) begin
        _tmp_900 <= _tmp_899;
      end 
      if(_mystream_stream_oready) begin
        _tmp_901 <= _tmp_900;
      end 
      if(_tmp_887) begin
        _mystream_sum_vec24_sink_mode <= 5'b1;
        _mystream_sum_vec24_sink_offset <= _tmp_893;
        _mystream_sum_vec24_sink_size <= _tmp_901;
        _mystream_sum_vec24_sink_stride <= 1;
      end 
      if(_tmp_887) begin
        _mystream_sum_vec24_sink_sel <= 89;
      end 
      if(_mystream_sink_start && _mystream_sum_vec24_sink_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_sum_vec24_sink_offset_buf <= _mystream_sum_vec24_sink_offset;
        _mystream_sum_vec24_sink_size_buf <= _mystream_sum_vec24_sink_size;
        _mystream_sum_vec24_sink_stride_buf <= _mystream_sum_vec24_sink_stride;
      end 
      if((_mystream_sum_vec24_sink_fsm_88 == 1) && _mystream_stream_oready) begin
        _mystream_sum_vec24_sink_waddr <= _mystream_sum_vec24_sink_offset_buf - _mystream_sum_vec24_sink_stride_buf;
        _mystream_sum_vec24_sink_count <= _mystream_sum_vec24_sink_size_buf;
      end 
      if((_mystream_sum_vec24_sink_fsm_88 == 2) && _mystream_stream_oready) begin
        _mystream_sum_vec24_sink_waddr <= _mystream_sum_vec24_sink_waddr + _mystream_sum_vec24_sink_stride_buf;
        _mystream_sum_vec24_sink_wdata <= mystream_sum_vec24_data;
        _mystream_sum_vec24_sink_wenable <= 1;
        _mystream_sum_vec24_sink_count <= _mystream_sum_vec24_sink_count - 1;
      end 
      if(_mystream_stream_oready) begin
        _tmp_903 <= _set_flag_902;
      end 
      if(_mystream_stream_oready) begin
        _tmp_904 <= _tmp_903;
      end 
      if(_mystream_stream_oready) begin
        _tmp_905 <= _tmp_904;
      end 
      if(_mystream_stream_oready) begin
        _tmp_906 <= _tmp_905;
      end 
      if(_mystream_stream_oready) begin
        _tmp_907 <= _tmp_906;
      end 
      if(_mystream_stream_oready) begin
        _tmp_908 <= _tmp_907;
      end 
      if(_mystream_stream_oready) begin
        _tmp_909 <= _th_comp_offset_4;
      end 
      if(_mystream_stream_oready) begin
        _tmp_910 <= _tmp_909;
      end 
      if(_mystream_stream_oready) begin
        _tmp_911 <= _tmp_910;
      end 
      if(_mystream_stream_oready) begin
        _tmp_912 <= _tmp_911;
      end 
      if(_mystream_stream_oready) begin
        _tmp_913 <= _tmp_912;
      end 
      if(_mystream_stream_oready) begin
        _tmp_914 <= _tmp_913;
      end 
      if(_mystream_stream_oready) begin
        _tmp_917 <= _tmp_916;
      end 
      if(_mystream_stream_oready) begin
        _tmp_918 <= _tmp_917;
      end 
      if(_mystream_stream_oready) begin
        _tmp_919 <= _tmp_918;
      end 
      if(_mystream_stream_oready) begin
        _tmp_920 <= _tmp_919;
      end 
      if(_mystream_stream_oready) begin
        _tmp_921 <= _tmp_920;
      end 
      if(_mystream_stream_oready) begin
        _tmp_922 <= _tmp_921;
      end 
      if(_tmp_908) begin
        _mystream_sum_vec25_sink_mode <= 5'b1;
        _mystream_sum_vec25_sink_offset <= _tmp_914;
        _mystream_sum_vec25_sink_size <= _tmp_922;
        _mystream_sum_vec25_sink_stride <= 1;
      end 
      if(_tmp_908) begin
        _mystream_sum_vec25_sink_sel <= 90;
      end 
      if(_mystream_sink_start && _mystream_sum_vec25_sink_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_sum_vec25_sink_offset_buf <= _mystream_sum_vec25_sink_offset;
        _mystream_sum_vec25_sink_size_buf <= _mystream_sum_vec25_sink_size;
        _mystream_sum_vec25_sink_stride_buf <= _mystream_sum_vec25_sink_stride;
      end 
      if((_mystream_sum_vec25_sink_fsm_89 == 1) && _mystream_stream_oready) begin
        _mystream_sum_vec25_sink_waddr <= _mystream_sum_vec25_sink_offset_buf - _mystream_sum_vec25_sink_stride_buf;
        _mystream_sum_vec25_sink_count <= _mystream_sum_vec25_sink_size_buf;
      end 
      if((_mystream_sum_vec25_sink_fsm_89 == 2) && _mystream_stream_oready) begin
        _mystream_sum_vec25_sink_waddr <= _mystream_sum_vec25_sink_waddr + _mystream_sum_vec25_sink_stride_buf;
        _mystream_sum_vec25_sink_wdata <= mystream_sum_vec25_data;
        _mystream_sum_vec25_sink_wenable <= 1;
        _mystream_sum_vec25_sink_count <= _mystream_sum_vec25_sink_count - 1;
      end 
      if(_mystream_stream_oready) begin
        _tmp_924 <= _set_flag_923;
      end 
      if(_mystream_stream_oready) begin
        _tmp_925 <= _tmp_924;
      end 
      if(_mystream_stream_oready) begin
        _tmp_926 <= _tmp_925;
      end 
      if(_mystream_stream_oready) begin
        _tmp_927 <= _tmp_926;
      end 
      if(_mystream_stream_oready) begin
        _tmp_928 <= _tmp_927;
      end 
      if(_mystream_stream_oready) begin
        _tmp_929 <= _tmp_928;
      end 
      if(_mystream_stream_oready) begin
        _tmp_930 <= _th_comp_offset_4;
      end 
      if(_mystream_stream_oready) begin
        _tmp_931 <= _tmp_930;
      end 
      if(_mystream_stream_oready) begin
        _tmp_932 <= _tmp_931;
      end 
      if(_mystream_stream_oready) begin
        _tmp_933 <= _tmp_932;
      end 
      if(_mystream_stream_oready) begin
        _tmp_934 <= _tmp_933;
      end 
      if(_mystream_stream_oready) begin
        _tmp_935 <= _tmp_934;
      end 
      if(_mystream_stream_oready) begin
        _tmp_938 <= _tmp_937;
      end 
      if(_mystream_stream_oready) begin
        _tmp_939 <= _tmp_938;
      end 
      if(_mystream_stream_oready) begin
        _tmp_940 <= _tmp_939;
      end 
      if(_mystream_stream_oready) begin
        _tmp_941 <= _tmp_940;
      end 
      if(_mystream_stream_oready) begin
        _tmp_942 <= _tmp_941;
      end 
      if(_mystream_stream_oready) begin
        _tmp_943 <= _tmp_942;
      end 
      if(_tmp_929) begin
        _mystream_sum_vec26_sink_mode <= 5'b1;
        _mystream_sum_vec26_sink_offset <= _tmp_935;
        _mystream_sum_vec26_sink_size <= _tmp_943;
        _mystream_sum_vec26_sink_stride <= 1;
      end 
      if(_tmp_929) begin
        _mystream_sum_vec26_sink_sel <= 91;
      end 
      if(_mystream_sink_start && _mystream_sum_vec26_sink_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_sum_vec26_sink_offset_buf <= _mystream_sum_vec26_sink_offset;
        _mystream_sum_vec26_sink_size_buf <= _mystream_sum_vec26_sink_size;
        _mystream_sum_vec26_sink_stride_buf <= _mystream_sum_vec26_sink_stride;
      end 
      if((_mystream_sum_vec26_sink_fsm_90 == 1) && _mystream_stream_oready) begin
        _mystream_sum_vec26_sink_waddr <= _mystream_sum_vec26_sink_offset_buf - _mystream_sum_vec26_sink_stride_buf;
        _mystream_sum_vec26_sink_count <= _mystream_sum_vec26_sink_size_buf;
      end 
      if((_mystream_sum_vec26_sink_fsm_90 == 2) && _mystream_stream_oready) begin
        _mystream_sum_vec26_sink_waddr <= _mystream_sum_vec26_sink_waddr + _mystream_sum_vec26_sink_stride_buf;
        _mystream_sum_vec26_sink_wdata <= mystream_sum_vec26_data;
        _mystream_sum_vec26_sink_wenable <= 1;
        _mystream_sum_vec26_sink_count <= _mystream_sum_vec26_sink_count - 1;
      end 
      if(_mystream_stream_oready) begin
        _tmp_945 <= _set_flag_944;
      end 
      if(_mystream_stream_oready) begin
        _tmp_946 <= _tmp_945;
      end 
      if(_mystream_stream_oready) begin
        _tmp_947 <= _tmp_946;
      end 
      if(_mystream_stream_oready) begin
        _tmp_948 <= _tmp_947;
      end 
      if(_mystream_stream_oready) begin
        _tmp_949 <= _tmp_948;
      end 
      if(_mystream_stream_oready) begin
        _tmp_950 <= _tmp_949;
      end 
      if(_mystream_stream_oready) begin
        _tmp_951 <= _th_comp_offset_4;
      end 
      if(_mystream_stream_oready) begin
        _tmp_952 <= _tmp_951;
      end 
      if(_mystream_stream_oready) begin
        _tmp_953 <= _tmp_952;
      end 
      if(_mystream_stream_oready) begin
        _tmp_954 <= _tmp_953;
      end 
      if(_mystream_stream_oready) begin
        _tmp_955 <= _tmp_954;
      end 
      if(_mystream_stream_oready) begin
        _tmp_956 <= _tmp_955;
      end 
      if(_mystream_stream_oready) begin
        _tmp_959 <= _tmp_958;
      end 
      if(_mystream_stream_oready) begin
        _tmp_960 <= _tmp_959;
      end 
      if(_mystream_stream_oready) begin
        _tmp_961 <= _tmp_960;
      end 
      if(_mystream_stream_oready) begin
        _tmp_962 <= _tmp_961;
      end 
      if(_mystream_stream_oready) begin
        _tmp_963 <= _tmp_962;
      end 
      if(_mystream_stream_oready) begin
        _tmp_964 <= _tmp_963;
      end 
      if(_tmp_950) begin
        _mystream_sum_vec27_sink_mode <= 5'b1;
        _mystream_sum_vec27_sink_offset <= _tmp_956;
        _mystream_sum_vec27_sink_size <= _tmp_964;
        _mystream_sum_vec27_sink_stride <= 1;
      end 
      if(_tmp_950) begin
        _mystream_sum_vec27_sink_sel <= 92;
      end 
      if(_mystream_sink_start && _mystream_sum_vec27_sink_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_sum_vec27_sink_offset_buf <= _mystream_sum_vec27_sink_offset;
        _mystream_sum_vec27_sink_size_buf <= _mystream_sum_vec27_sink_size;
        _mystream_sum_vec27_sink_stride_buf <= _mystream_sum_vec27_sink_stride;
      end 
      if((_mystream_sum_vec27_sink_fsm_91 == 1) && _mystream_stream_oready) begin
        _mystream_sum_vec27_sink_waddr <= _mystream_sum_vec27_sink_offset_buf - _mystream_sum_vec27_sink_stride_buf;
        _mystream_sum_vec27_sink_count <= _mystream_sum_vec27_sink_size_buf;
      end 
      if((_mystream_sum_vec27_sink_fsm_91 == 2) && _mystream_stream_oready) begin
        _mystream_sum_vec27_sink_waddr <= _mystream_sum_vec27_sink_waddr + _mystream_sum_vec27_sink_stride_buf;
        _mystream_sum_vec27_sink_wdata <= mystream_sum_vec27_data;
        _mystream_sum_vec27_sink_wenable <= 1;
        _mystream_sum_vec27_sink_count <= _mystream_sum_vec27_sink_count - 1;
      end 
      if(_mystream_stream_oready) begin
        _tmp_966 <= _set_flag_965;
      end 
      if(_mystream_stream_oready) begin
        _tmp_967 <= _tmp_966;
      end 
      if(_mystream_stream_oready) begin
        _tmp_968 <= _tmp_967;
      end 
      if(_mystream_stream_oready) begin
        _tmp_969 <= _tmp_968;
      end 
      if(_mystream_stream_oready) begin
        _tmp_970 <= _tmp_969;
      end 
      if(_mystream_stream_oready) begin
        _tmp_971 <= _tmp_970;
      end 
      if(_mystream_stream_oready) begin
        _tmp_972 <= _th_comp_offset_4;
      end 
      if(_mystream_stream_oready) begin
        _tmp_973 <= _tmp_972;
      end 
      if(_mystream_stream_oready) begin
        _tmp_974 <= _tmp_973;
      end 
      if(_mystream_stream_oready) begin
        _tmp_975 <= _tmp_974;
      end 
      if(_mystream_stream_oready) begin
        _tmp_976 <= _tmp_975;
      end 
      if(_mystream_stream_oready) begin
        _tmp_977 <= _tmp_976;
      end 
      if(_mystream_stream_oready) begin
        _tmp_980 <= _tmp_979;
      end 
      if(_mystream_stream_oready) begin
        _tmp_981 <= _tmp_980;
      end 
      if(_mystream_stream_oready) begin
        _tmp_982 <= _tmp_981;
      end 
      if(_mystream_stream_oready) begin
        _tmp_983 <= _tmp_982;
      end 
      if(_mystream_stream_oready) begin
        _tmp_984 <= _tmp_983;
      end 
      if(_mystream_stream_oready) begin
        _tmp_985 <= _tmp_984;
      end 
      if(_tmp_971) begin
        _mystream_sum_vec28_sink_mode <= 5'b1;
        _mystream_sum_vec28_sink_offset <= _tmp_977;
        _mystream_sum_vec28_sink_size <= _tmp_985;
        _mystream_sum_vec28_sink_stride <= 1;
      end 
      if(_tmp_971) begin
        _mystream_sum_vec28_sink_sel <= 93;
      end 
      if(_mystream_sink_start && _mystream_sum_vec28_sink_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_sum_vec28_sink_offset_buf <= _mystream_sum_vec28_sink_offset;
        _mystream_sum_vec28_sink_size_buf <= _mystream_sum_vec28_sink_size;
        _mystream_sum_vec28_sink_stride_buf <= _mystream_sum_vec28_sink_stride;
      end 
      if((_mystream_sum_vec28_sink_fsm_92 == 1) && _mystream_stream_oready) begin
        _mystream_sum_vec28_sink_waddr <= _mystream_sum_vec28_sink_offset_buf - _mystream_sum_vec28_sink_stride_buf;
        _mystream_sum_vec28_sink_count <= _mystream_sum_vec28_sink_size_buf;
      end 
      if((_mystream_sum_vec28_sink_fsm_92 == 2) && _mystream_stream_oready) begin
        _mystream_sum_vec28_sink_waddr <= _mystream_sum_vec28_sink_waddr + _mystream_sum_vec28_sink_stride_buf;
        _mystream_sum_vec28_sink_wdata <= mystream_sum_vec28_data;
        _mystream_sum_vec28_sink_wenable <= 1;
        _mystream_sum_vec28_sink_count <= _mystream_sum_vec28_sink_count - 1;
      end 
      if(_mystream_stream_oready) begin
        _tmp_987 <= _set_flag_986;
      end 
      if(_mystream_stream_oready) begin
        _tmp_988 <= _tmp_987;
      end 
      if(_mystream_stream_oready) begin
        _tmp_989 <= _tmp_988;
      end 
      if(_mystream_stream_oready) begin
        _tmp_990 <= _tmp_989;
      end 
      if(_mystream_stream_oready) begin
        _tmp_991 <= _tmp_990;
      end 
      if(_mystream_stream_oready) begin
        _tmp_992 <= _tmp_991;
      end 
      if(_mystream_stream_oready) begin
        _tmp_993 <= _th_comp_offset_4;
      end 
      if(_mystream_stream_oready) begin
        _tmp_994 <= _tmp_993;
      end 
      if(_mystream_stream_oready) begin
        _tmp_995 <= _tmp_994;
      end 
      if(_mystream_stream_oready) begin
        _tmp_996 <= _tmp_995;
      end 
      if(_mystream_stream_oready) begin
        _tmp_997 <= _tmp_996;
      end 
      if(_mystream_stream_oready) begin
        _tmp_998 <= _tmp_997;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1001 <= _tmp_1000;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1002 <= _tmp_1001;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1003 <= _tmp_1002;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1004 <= _tmp_1003;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1005 <= _tmp_1004;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1006 <= _tmp_1005;
      end 
      if(_tmp_992) begin
        _mystream_sum_vec29_sink_mode <= 5'b1;
        _mystream_sum_vec29_sink_offset <= _tmp_998;
        _mystream_sum_vec29_sink_size <= _tmp_1006;
        _mystream_sum_vec29_sink_stride <= 1;
      end 
      if(_tmp_992) begin
        _mystream_sum_vec29_sink_sel <= 94;
      end 
      if(_mystream_sink_start && _mystream_sum_vec29_sink_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_sum_vec29_sink_offset_buf <= _mystream_sum_vec29_sink_offset;
        _mystream_sum_vec29_sink_size_buf <= _mystream_sum_vec29_sink_size;
        _mystream_sum_vec29_sink_stride_buf <= _mystream_sum_vec29_sink_stride;
      end 
      if((_mystream_sum_vec29_sink_fsm_93 == 1) && _mystream_stream_oready) begin
        _mystream_sum_vec29_sink_waddr <= _mystream_sum_vec29_sink_offset_buf - _mystream_sum_vec29_sink_stride_buf;
        _mystream_sum_vec29_sink_count <= _mystream_sum_vec29_sink_size_buf;
      end 
      if((_mystream_sum_vec29_sink_fsm_93 == 2) && _mystream_stream_oready) begin
        _mystream_sum_vec29_sink_waddr <= _mystream_sum_vec29_sink_waddr + _mystream_sum_vec29_sink_stride_buf;
        _mystream_sum_vec29_sink_wdata <= mystream_sum_vec29_data;
        _mystream_sum_vec29_sink_wenable <= 1;
        _mystream_sum_vec29_sink_count <= _mystream_sum_vec29_sink_count - 1;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1008 <= _set_flag_1007;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1009 <= _tmp_1008;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1010 <= _tmp_1009;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1011 <= _tmp_1010;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1012 <= _tmp_1011;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1013 <= _tmp_1012;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1014 <= _th_comp_offset_4;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1015 <= _tmp_1014;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1016 <= _tmp_1015;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1017 <= _tmp_1016;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1018 <= _tmp_1017;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1019 <= _tmp_1018;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1022 <= _tmp_1021;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1023 <= _tmp_1022;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1024 <= _tmp_1023;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1025 <= _tmp_1024;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1026 <= _tmp_1025;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1027 <= _tmp_1026;
      end 
      if(_tmp_1013) begin
        _mystream_sum_vec30_sink_mode <= 5'b1;
        _mystream_sum_vec30_sink_offset <= _tmp_1019;
        _mystream_sum_vec30_sink_size <= _tmp_1027;
        _mystream_sum_vec30_sink_stride <= 1;
      end 
      if(_tmp_1013) begin
        _mystream_sum_vec30_sink_sel <= 95;
      end 
      if(_mystream_sink_start && _mystream_sum_vec30_sink_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_sum_vec30_sink_offset_buf <= _mystream_sum_vec30_sink_offset;
        _mystream_sum_vec30_sink_size_buf <= _mystream_sum_vec30_sink_size;
        _mystream_sum_vec30_sink_stride_buf <= _mystream_sum_vec30_sink_stride;
      end 
      if((_mystream_sum_vec30_sink_fsm_94 == 1) && _mystream_stream_oready) begin
        _mystream_sum_vec30_sink_waddr <= _mystream_sum_vec30_sink_offset_buf - _mystream_sum_vec30_sink_stride_buf;
        _mystream_sum_vec30_sink_count <= _mystream_sum_vec30_sink_size_buf;
      end 
      if((_mystream_sum_vec30_sink_fsm_94 == 2) && _mystream_stream_oready) begin
        _mystream_sum_vec30_sink_waddr <= _mystream_sum_vec30_sink_waddr + _mystream_sum_vec30_sink_stride_buf;
        _mystream_sum_vec30_sink_wdata <= mystream_sum_vec30_data;
        _mystream_sum_vec30_sink_wenable <= 1;
        _mystream_sum_vec30_sink_count <= _mystream_sum_vec30_sink_count - 1;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1029 <= _set_flag_1028;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1030 <= _tmp_1029;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1031 <= _tmp_1030;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1032 <= _tmp_1031;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1033 <= _tmp_1032;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1034 <= _tmp_1033;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1035 <= _th_comp_offset_4;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1036 <= _tmp_1035;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1037 <= _tmp_1036;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1038 <= _tmp_1037;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1039 <= _tmp_1038;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1040 <= _tmp_1039;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1043 <= _tmp_1042;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1044 <= _tmp_1043;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1045 <= _tmp_1044;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1046 <= _tmp_1045;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1047 <= _tmp_1046;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1048 <= _tmp_1047;
      end 
      if(_tmp_1034) begin
        _mystream_sum_vec31_sink_mode <= 5'b1;
        _mystream_sum_vec31_sink_offset <= _tmp_1040;
        _mystream_sum_vec31_sink_size <= _tmp_1048;
        _mystream_sum_vec31_sink_stride <= 1;
      end 
      if(_tmp_1034) begin
        _mystream_sum_vec31_sink_sel <= 96;
      end 
      if(_mystream_sink_start && _mystream_sum_vec31_sink_mode & 5'b1 && _mystream_stream_oready) begin
        _mystream_sum_vec31_sink_offset_buf <= _mystream_sum_vec31_sink_offset;
        _mystream_sum_vec31_sink_size_buf <= _mystream_sum_vec31_sink_size;
        _mystream_sum_vec31_sink_stride_buf <= _mystream_sum_vec31_sink_stride;
      end 
      if((_mystream_sum_vec31_sink_fsm_95 == 1) && _mystream_stream_oready) begin
        _mystream_sum_vec31_sink_waddr <= _mystream_sum_vec31_sink_offset_buf - _mystream_sum_vec31_sink_stride_buf;
        _mystream_sum_vec31_sink_count <= _mystream_sum_vec31_sink_size_buf;
      end 
      if((_mystream_sum_vec31_sink_fsm_95 == 2) && _mystream_stream_oready) begin
        _mystream_sum_vec31_sink_waddr <= _mystream_sum_vec31_sink_waddr + _mystream_sum_vec31_sink_stride_buf;
        _mystream_sum_vec31_sink_wdata <= mystream_sum_vec31_data;
        _mystream_sum_vec31_sink_wenable <= 1;
        _mystream_sum_vec31_sink_count <= _mystream_sum_vec31_sink_count - 1;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1050 <= _mystream_source_start;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1051 <= _tmp_1050;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1052 <= _tmp_1051;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1053 <= _mystream_source_start;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1054 <= _tmp_1053;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1055 <= _tmp_1054;
      end 
      if(_mystream_stream_oready && _tmp_1055) begin
        __variable_wdata_130 <= 1;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1056 <= _mystream_source_start;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1057 <= _tmp_1056;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1058 <= _tmp_1057;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1059 <= _tmp_1058;
      end 
      if(_mystream_stream_oready && _tmp_1059) begin
        __variable_wdata_130 <= 0;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1062 <= _tmp_1061;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1065 <= _tmp_1064;
      end 
      if(_mystream_stream_oready && _tmp_1065) begin
        __variable_wdata_130 <= 1;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1066 <= _mystream_source_start;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1067 <= _tmp_1066;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1068 <= _tmp_1067;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1069 <= _tmp_1068;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1070 <= _tmp_1069;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1071 <= _tmp_1070;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1072 <= _mystream_source_stop;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1073 <= _tmp_1072;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1074 <= _tmp_1073;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1075 <= _tmp_1074;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1076 <= _tmp_1075;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1077 <= _tmp_1076;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1078 <= _mystream_source_busy;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1079 <= _tmp_1078;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1080 <= _tmp_1079;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1081 <= _tmp_1080;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1082 <= _tmp_1081;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1083 <= _tmp_1082;
      end 
      if(_mystream_stream_oready) begin
        _tmp_1084 <= _mystream_sink_busy;
      end 
      if(!_mystream_sink_busy && _tmp_1084) begin
        _mystream_busy_reg <= 0;
      end 
      if(_mystream_source_busy) begin
        _mystream_busy_reg <= 1;
      end 
    end
  end

  localparam _mystream_fsm_1 = 1;
  localparam _mystream_fsm_2 = 2;
  localparam _mystream_fsm_3 = 3;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_fsm <= _mystream_fsm_init;
      _mystream_source_start <= 0;
      _mystream_source_busy <= 0;
      _mystream_stream_ivalid <= 0;
    end else begin
      if(_mystream_stream_oready && _tmp_1052) begin
        _mystream_stream_ivalid <= 1;
      end 
      if(_mystream_stream_oready && _tmp_1062) begin
        _mystream_stream_ivalid <= 0;
      end 
      case(_mystream_fsm)
        _mystream_fsm_init: begin
          if(_mystream_run_flag) begin
            _mystream_source_start <= 1;
          end 
          if(_mystream_run_flag) begin
            _mystream_fsm <= _mystream_fsm_1;
          end 
        end
        _mystream_fsm_1: begin
          if(_mystream_source_start && _mystream_stream_oready) begin
            _mystream_source_start <= 0;
            _mystream_source_busy <= 1;
          end 
          if(_mystream_source_start && _mystream_stream_oready) begin
            _mystream_fsm <= _mystream_fsm_2;
          end 
        end
        _mystream_fsm_2: begin
          if(_mystream_stream_oready) begin
            _mystream_fsm <= _mystream_fsm_3;
          end 
        end
        _mystream_fsm_3: begin
          if(_mystream_stream_oready && (_mystream_a0_idle && _mystream_a1_idle && _mystream_a10_idle && _mystream_a11_idle && _mystream_a12_idle && _mystream_a13_idle && _mystream_a14_idle && _mystream_a15_idle && _mystream_a16_idle && _mystream_a17_idle && _mystream_a18_idle && _mystream_a19_idle && _mystream_a2_idle && _mystream_a20_idle && _mystream_a21_idle && _mystream_a22_idle && _mystream_a23_idle && _mystream_a24_idle && _mystream_a25_idle && _mystream_a26_idle && _mystream_a27_idle && _mystream_a28_idle && _mystream_a29_idle && _mystream_a3_idle && _mystream_a30_idle && _mystream_a31_idle && _mystream_a4_idle && _mystream_a5_idle && _mystream_a6_idle && _mystream_a7_idle && _mystream_a8_idle && _mystream_a9_idle && _mystream_b0_idle && _mystream_b1_idle && _mystream_b10_idle && _mystream_b11_idle && _mystream_b12_idle && _mystream_b13_idle && _mystream_b14_idle && _mystream_b15_idle && _mystream_b16_idle && _mystream_b17_idle && _mystream_b18_idle && _mystream_b19_idle && _mystream_b2_idle && _mystream_b20_idle && _mystream_b21_idle && _mystream_b22_idle && _mystream_b23_idle && _mystream_b24_idle && _mystream_b25_idle && _mystream_b26_idle && _mystream_b27_idle && _mystream_b28_idle && _mystream_b29_idle && _mystream_b3_idle && _mystream_b30_idle && _mystream_b31_idle && _mystream_b4_idle && _mystream_b5_idle && _mystream_b6_idle && _mystream_b7_idle && _mystream_b8_idle && _mystream_b9_idle && _mystream_bias0_idle && _mystream_bias1_idle && _mystream_bias10_idle && _mystream_bias11_idle && _mystream_bias12_idle && _mystream_bias13_idle && _mystream_bias14_idle && _mystream_bias15_idle && _mystream_bias16_idle && _mystream_bias17_idle && _mystream_bias18_idle && _mystream_bias19_idle && _mystream_bias2_idle && _mystream_bias20_idle && _mystream_bias21_idle && _mystream_bias22_idle && _mystream_bias23_idle && _mystream_bias24_idle && _mystream_bias25_idle && _mystream_bias26_idle && _mystream_bias27_idle && _mystream_bias28_idle && _mystream_bias29_idle && _mystream_bias3_idle && _mystream_bias30_idle && _mystream_bias31_idle && _mystream_bias4_idle && _mystream_bias5_idle && _mystream_bias6_idle && _mystream_bias7_idle && _mystream_bias8_idle && _mystream_bias9_idle && (_mystream_fsm == 3))) begin
            _mystream_source_busy <= 0;
          end 
          if(_mystream_stream_oready && (_mystream_a0_idle && _mystream_a1_idle && _mystream_a10_idle && _mystream_a11_idle && _mystream_a12_idle && _mystream_a13_idle && _mystream_a14_idle && _mystream_a15_idle && _mystream_a16_idle && _mystream_a17_idle && _mystream_a18_idle && _mystream_a19_idle && _mystream_a2_idle && _mystream_a20_idle && _mystream_a21_idle && _mystream_a22_idle && _mystream_a23_idle && _mystream_a24_idle && _mystream_a25_idle && _mystream_a26_idle && _mystream_a27_idle && _mystream_a28_idle && _mystream_a29_idle && _mystream_a3_idle && _mystream_a30_idle && _mystream_a31_idle && _mystream_a4_idle && _mystream_a5_idle && _mystream_a6_idle && _mystream_a7_idle && _mystream_a8_idle && _mystream_a9_idle && _mystream_b0_idle && _mystream_b1_idle && _mystream_b10_idle && _mystream_b11_idle && _mystream_b12_idle && _mystream_b13_idle && _mystream_b14_idle && _mystream_b15_idle && _mystream_b16_idle && _mystream_b17_idle && _mystream_b18_idle && _mystream_b19_idle && _mystream_b2_idle && _mystream_b20_idle && _mystream_b21_idle && _mystream_b22_idle && _mystream_b23_idle && _mystream_b24_idle && _mystream_b25_idle && _mystream_b26_idle && _mystream_b27_idle && _mystream_b28_idle && _mystream_b29_idle && _mystream_b3_idle && _mystream_b30_idle && _mystream_b31_idle && _mystream_b4_idle && _mystream_b5_idle && _mystream_b6_idle && _mystream_b7_idle && _mystream_b8_idle && _mystream_b9_idle && _mystream_bias0_idle && _mystream_bias1_idle && _mystream_bias10_idle && _mystream_bias11_idle && _mystream_bias12_idle && _mystream_bias13_idle && _mystream_bias14_idle && _mystream_bias15_idle && _mystream_bias16_idle && _mystream_bias17_idle && _mystream_bias18_idle && _mystream_bias19_idle && _mystream_bias2_idle && _mystream_bias20_idle && _mystream_bias21_idle && _mystream_bias22_idle && _mystream_bias23_idle && _mystream_bias24_idle && _mystream_bias25_idle && _mystream_bias26_idle && _mystream_bias27_idle && _mystream_bias28_idle && _mystream_bias29_idle && _mystream_bias3_idle && _mystream_bias30_idle && _mystream_bias31_idle && _mystream_bias4_idle && _mystream_bias5_idle && _mystream_bias6_idle && _mystream_bias7_idle && _mystream_bias8_idle && _mystream_bias9_idle && (_mystream_fsm == 3)) && _mystream_run_flag) begin
            _mystream_source_start <= 1;
          end 
          if(_mystream_stream_oready && (_mystream_a0_idle && _mystream_a1_idle && _mystream_a10_idle && _mystream_a11_idle && _mystream_a12_idle && _mystream_a13_idle && _mystream_a14_idle && _mystream_a15_idle && _mystream_a16_idle && _mystream_a17_idle && _mystream_a18_idle && _mystream_a19_idle && _mystream_a2_idle && _mystream_a20_idle && _mystream_a21_idle && _mystream_a22_idle && _mystream_a23_idle && _mystream_a24_idle && _mystream_a25_idle && _mystream_a26_idle && _mystream_a27_idle && _mystream_a28_idle && _mystream_a29_idle && _mystream_a3_idle && _mystream_a30_idle && _mystream_a31_idle && _mystream_a4_idle && _mystream_a5_idle && _mystream_a6_idle && _mystream_a7_idle && _mystream_a8_idle && _mystream_a9_idle && _mystream_b0_idle && _mystream_b1_idle && _mystream_b10_idle && _mystream_b11_idle && _mystream_b12_idle && _mystream_b13_idle && _mystream_b14_idle && _mystream_b15_idle && _mystream_b16_idle && _mystream_b17_idle && _mystream_b18_idle && _mystream_b19_idle && _mystream_b2_idle && _mystream_b20_idle && _mystream_b21_idle && _mystream_b22_idle && _mystream_b23_idle && _mystream_b24_idle && _mystream_b25_idle && _mystream_b26_idle && _mystream_b27_idle && _mystream_b28_idle && _mystream_b29_idle && _mystream_b3_idle && _mystream_b30_idle && _mystream_b31_idle && _mystream_b4_idle && _mystream_b5_idle && _mystream_b6_idle && _mystream_b7_idle && _mystream_b8_idle && _mystream_b9_idle && _mystream_bias0_idle && _mystream_bias1_idle && _mystream_bias10_idle && _mystream_bias11_idle && _mystream_bias12_idle && _mystream_bias13_idle && _mystream_bias14_idle && _mystream_bias15_idle && _mystream_bias16_idle && _mystream_bias17_idle && _mystream_bias18_idle && _mystream_bias19_idle && _mystream_bias2_idle && _mystream_bias20_idle && _mystream_bias21_idle && _mystream_bias22_idle && _mystream_bias23_idle && _mystream_bias24_idle && _mystream_bias25_idle && _mystream_bias26_idle && _mystream_bias27_idle && _mystream_bias28_idle && _mystream_bias29_idle && _mystream_bias3_idle && _mystream_bias30_idle && _mystream_bias31_idle && _mystream_bias4_idle && _mystream_bias5_idle && _mystream_bias6_idle && _mystream_bias7_idle && _mystream_bias8_idle && _mystream_bias9_idle && (_mystream_fsm == 3))) begin
            _mystream_fsm <= _mystream_fsm_init;
          end 
          if(_mystream_stream_oready && (_mystream_a0_idle && _mystream_a1_idle && _mystream_a10_idle && _mystream_a11_idle && _mystream_a12_idle && _mystream_a13_idle && _mystream_a14_idle && _mystream_a15_idle && _mystream_a16_idle && _mystream_a17_idle && _mystream_a18_idle && _mystream_a19_idle && _mystream_a2_idle && _mystream_a20_idle && _mystream_a21_idle && _mystream_a22_idle && _mystream_a23_idle && _mystream_a24_idle && _mystream_a25_idle && _mystream_a26_idle && _mystream_a27_idle && _mystream_a28_idle && _mystream_a29_idle && _mystream_a3_idle && _mystream_a30_idle && _mystream_a31_idle && _mystream_a4_idle && _mystream_a5_idle && _mystream_a6_idle && _mystream_a7_idle && _mystream_a8_idle && _mystream_a9_idle && _mystream_b0_idle && _mystream_b1_idle && _mystream_b10_idle && _mystream_b11_idle && _mystream_b12_idle && _mystream_b13_idle && _mystream_b14_idle && _mystream_b15_idle && _mystream_b16_idle && _mystream_b17_idle && _mystream_b18_idle && _mystream_b19_idle && _mystream_b2_idle && _mystream_b20_idle && _mystream_b21_idle && _mystream_b22_idle && _mystream_b23_idle && _mystream_b24_idle && _mystream_b25_idle && _mystream_b26_idle && _mystream_b27_idle && _mystream_b28_idle && _mystream_b29_idle && _mystream_b3_idle && _mystream_b30_idle && _mystream_b31_idle && _mystream_b4_idle && _mystream_b5_idle && _mystream_b6_idle && _mystream_b7_idle && _mystream_b8_idle && _mystream_b9_idle && _mystream_bias0_idle && _mystream_bias1_idle && _mystream_bias10_idle && _mystream_bias11_idle && _mystream_bias12_idle && _mystream_bias13_idle && _mystream_bias14_idle && _mystream_bias15_idle && _mystream_bias16_idle && _mystream_bias17_idle && _mystream_bias18_idle && _mystream_bias19_idle && _mystream_bias2_idle && _mystream_bias20_idle && _mystream_bias21_idle && _mystream_bias22_idle && _mystream_bias23_idle && _mystream_bias24_idle && _mystream_bias25_idle && _mystream_bias26_idle && _mystream_bias27_idle && _mystream_bias28_idle && _mystream_bias29_idle && _mystream_bias3_idle && _mystream_bias30_idle && _mystream_bias31_idle && _mystream_bias4_idle && _mystream_bias5_idle && _mystream_bias6_idle && _mystream_bias7_idle && _mystream_bias8_idle && _mystream_bias9_idle && (_mystream_fsm == 3)) && _mystream_run_flag) begin
            _mystream_fsm <= _mystream_fsm_1;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      counter <= 0;
    end else begin
      counter <= counter + 1;
    end
  end

  localparam th_comp_1 = 1;
  localparam th_comp_2 = 2;
  localparam th_comp_3 = 3;
  localparam th_comp_4 = 4;
  localparam th_comp_5 = 5;
  localparam th_comp_6 = 6;
  localparam th_comp_7 = 7;
  localparam th_comp_8 = 8;
  localparam th_comp_9 = 9;
  localparam th_comp_10 = 10;
  localparam th_comp_11 = 11;
  localparam th_comp_12 = 12;
  localparam th_comp_13 = 13;
  localparam th_comp_14 = 14;
  localparam th_comp_15 = 15;
  localparam th_comp_16 = 16;
  localparam th_comp_17 = 17;
  localparam th_comp_18 = 18;
  localparam th_comp_19 = 19;
  localparam th_comp_20 = 20;
  localparam th_comp_21 = 21;
  localparam th_comp_22 = 22;
  localparam th_comp_23 = 23;
  localparam th_comp_24 = 24;
  localparam th_comp_25 = 25;
  localparam th_comp_26 = 26;
  localparam th_comp_27 = 27;
  localparam th_comp_28 = 28;
  localparam th_comp_29 = 29;
  localparam th_comp_30 = 30;
  localparam th_comp_31 = 31;
  localparam th_comp_32 = 32;
  localparam th_comp_33 = 33;
  localparam th_comp_34 = 34;
  localparam th_comp_35 = 35;
  localparam th_comp_36 = 36;
  localparam th_comp_37 = 37;
  localparam th_comp_38 = 38;
  localparam th_comp_39 = 39;
  localparam th_comp_40 = 40;
  localparam th_comp_41 = 41;
  localparam th_comp_42 = 42;
  localparam th_comp_43 = 43;
  localparam th_comp_44 = 44;
  localparam th_comp_45 = 45;
  localparam th_comp_46 = 46;
  localparam th_comp_47 = 47;
  localparam th_comp_48 = 48;
  localparam th_comp_49 = 49;
  localparam th_comp_50 = 50;
  localparam th_comp_51 = 51;
  localparam th_comp_52 = 52;
  localparam th_comp_53 = 53;
  localparam th_comp_54 = 54;
  localparam th_comp_55 = 55;
  localparam th_comp_56 = 56;
  localparam th_comp_57 = 57;
  localparam th_comp_58 = 58;
  localparam th_comp_59 = 59;
  localparam th_comp_60 = 60;
  localparam th_comp_61 = 61;
  localparam th_comp_62 = 62;
  localparam th_comp_63 = 63;
  localparam th_comp_64 = 64;
  localparam th_comp_65 = 65;
  localparam th_comp_66 = 66;
  localparam th_comp_67 = 67;
  localparam th_comp_68 = 68;
  localparam th_comp_69 = 69;
  localparam th_comp_70 = 70;
  localparam th_comp_71 = 71;
  localparam th_comp_72 = 72;
  localparam th_comp_73 = 73;
  localparam th_comp_74 = 74;
  localparam th_comp_75 = 75;
  localparam th_comp_76 = 76;
  localparam th_comp_77 = 77;
  localparam th_comp_78 = 78;
  localparam th_comp_79 = 79;
  localparam th_comp_80 = 80;
  localparam th_comp_81 = 81;
  localparam th_comp_82 = 82;
  localparam th_comp_83 = 83;
  localparam th_comp_84 = 84;
  localparam th_comp_85 = 85;
  localparam th_comp_86 = 86;
  localparam th_comp_87 = 87;
  localparam th_comp_88 = 88;
  localparam th_comp_89 = 89;
  localparam th_comp_90 = 90;
  localparam th_comp_91 = 91;
  localparam th_comp_92 = 92;
  localparam th_comp_93 = 93;
  localparam th_comp_94 = 94;
  localparam th_comp_95 = 95;
  localparam th_comp_96 = 96;
  localparam th_comp_97 = 97;
  localparam th_comp_98 = 98;
  localparam th_comp_99 = 99;
  localparam th_comp_100 = 100;
  localparam th_comp_101 = 101;
  localparam th_comp_102 = 102;
  localparam th_comp_103 = 103;
  localparam th_comp_104 = 104;
  localparam th_comp_105 = 105;
  localparam th_comp_106 = 106;
  localparam th_comp_107 = 107;
  localparam th_comp_108 = 108;
  localparam th_comp_109 = 109;
  localparam th_comp_110 = 110;
  localparam th_comp_111 = 111;
  localparam th_comp_112 = 112;
  localparam th_comp_113 = 113;
  localparam th_comp_114 = 114;
  localparam th_comp_115 = 115;
  localparam th_comp_116 = 116;
  localparam th_comp_117 = 117;
  localparam th_comp_118 = 118;
  localparam th_comp_119 = 119;
  localparam th_comp_120 = 120;
  localparam th_comp_121 = 121;
  localparam th_comp_122 = 122;
  localparam th_comp_123 = 123;
  localparam th_comp_124 = 124;
  localparam th_comp_125 = 125;
  localparam th_comp_126 = 126;

  always @(posedge CLK) begin
    if(RST) begin
      th_comp <= th_comp_init;
      _th_comp_size_0 <= 0;
      _th_comp_offset_b_1 <= 0;
      _th_comp_offset_2 <= 0;
      _th_comp_size_3 <= 0;
      _th_comp_offset_4 <= 0;
      _th_comp_start_time_5 <= 0;
      _th_comp_end_time_6 <= 0;
      _th_comp_exec_time_7 <= 0;
      _th_comp_size_8 <= 0;
      _th_comp_offset_9 <= 0;
      _th_comp_sum_10 <= 0;
      _th_comp_i_11 <= 0;
      read_rdata_1099 <= 0;
      _th_comp_a_12 <= 0;
      read_rdata_1102 <= 0;
      _th_comp_b_13 <= 0;
      _th_comp_size_14 <= 0;
      _th_comp_offset_stream_15 <= 0;
      _th_comp_offset_seq_16 <= 0;
      _th_comp_all_ok_17 <= 0;
      _th_comp_i_18 <= 0;
      read_rdata_1285 <= 0;
      _th_comp_st_19 <= 0;
      read_rdata_1354 <= 0;
      _th_comp_sq_20 <= 0;
    end else begin
      case(th_comp)
        th_comp_init: begin
          _th_comp_size_0 <= 1024;
          th_comp <= th_comp_1;
        end
        th_comp_1: begin
          _th_comp_offset_b_1 <= _th_comp_size_0 << 2;
          th_comp <= th_comp_2;
        end
        th_comp_2: begin
          _th_comp_size_0 <= _th_comp_size_0 >>> 1;
          th_comp <= th_comp_3;
        end
        th_comp_3: begin
          _th_comp_offset_2 <= 0;
          th_comp <= th_comp_4;
        end
        th_comp_4: begin
          if(_myaxi_read_req_idle) begin
            th_comp <= th_comp_5;
          end 
        end
        th_comp_5: begin
          if(_myaxi_read_idle) begin
            th_comp <= th_comp_6;
          end 
        end
        th_comp_6: begin
          if(_myaxi_read_req_idle) begin
            th_comp <= th_comp_7;
          end 
        end
        th_comp_7: begin
          if(_myaxi_read_idle) begin
            th_comp <= th_comp_8;
          end 
        end
        th_comp_8: begin
          _th_comp_size_3 <= _th_comp_size_0;
          _th_comp_offset_4 <= _th_comp_offset_2;
          th_comp <= th_comp_9;
        end
        th_comp_9: begin
          _th_comp_start_time_5 <= counter;
          th_comp <= th_comp_10;
        end
        th_comp_10: begin
          th_comp <= th_comp_11;
        end
        th_comp_11: begin
          th_comp <= th_comp_12;
        end
        th_comp_12: begin
          _th_comp_end_time_6 <= counter;
          th_comp <= th_comp_13;
        end
        th_comp_13: begin
          $display("# para = %d, exec_time = %d", 32, (_th_comp_end_time_6 - _th_comp_start_time_5));
          th_comp <= th_comp_14;
        end
        th_comp_14: begin
          th_comp <= th_comp_15;
        end
        th_comp_15: begin
          th_comp <= th_comp_16;
        end
        th_comp_16: begin
          th_comp <= th_comp_17;
        end
        th_comp_17: begin
          th_comp <= th_comp_18;
        end
        th_comp_18: begin
          th_comp <= th_comp_19;
        end
        th_comp_19: begin
          th_comp <= th_comp_20;
        end
        th_comp_20: begin
          th_comp <= th_comp_21;
        end
        th_comp_21: begin
          th_comp <= th_comp_22;
        end
        th_comp_22: begin
          th_comp <= th_comp_23;
        end
        th_comp_23: begin
          th_comp <= th_comp_24;
        end
        th_comp_24: begin
          th_comp <= th_comp_25;
        end
        th_comp_25: begin
          th_comp <= th_comp_26;
        end
        th_comp_26: begin
          th_comp <= th_comp_27;
        end
        th_comp_27: begin
          th_comp <= th_comp_28;
        end
        th_comp_28: begin
          th_comp <= th_comp_29;
        end
        th_comp_29: begin
          th_comp <= th_comp_30;
        end
        th_comp_30: begin
          th_comp <= th_comp_31;
        end
        th_comp_31: begin
          th_comp <= th_comp_32;
        end
        th_comp_32: begin
          th_comp <= th_comp_33;
        end
        th_comp_33: begin
          th_comp <= th_comp_34;
        end
        th_comp_34: begin
          th_comp <= th_comp_35;
        end
        th_comp_35: begin
          th_comp <= th_comp_36;
        end
        th_comp_36: begin
          th_comp <= th_comp_37;
        end
        th_comp_37: begin
          th_comp <= th_comp_38;
        end
        th_comp_38: begin
          th_comp <= th_comp_39;
        end
        th_comp_39: begin
          th_comp <= th_comp_40;
        end
        th_comp_40: begin
          th_comp <= th_comp_41;
        end
        th_comp_41: begin
          th_comp <= th_comp_42;
        end
        th_comp_42: begin
          th_comp <= th_comp_43;
        end
        th_comp_43: begin
          th_comp <= th_comp_44;
        end
        th_comp_44: begin
          th_comp <= th_comp_45;
        end
        th_comp_45: begin
          th_comp <= th_comp_46;
        end
        th_comp_46: begin
          _th_comp_end_time_6 <= counter;
          th_comp <= th_comp_47;
        end
        th_comp_47: begin
          $display("# para = %d, exec1_time = %d", 32, (_th_comp_end_time_6 - _th_comp_start_time_5));
          th_comp <= th_comp_48;
        end
        th_comp_48: begin
          th_comp <= th_comp_49;
        end
        th_comp_49: begin
          th_comp <= th_comp_50;
        end
        th_comp_50: begin
          th_comp <= th_comp_51;
        end
        th_comp_51: begin
          th_comp <= th_comp_52;
        end
        th_comp_52: begin
          th_comp <= th_comp_53;
        end
        th_comp_53: begin
          th_comp <= th_comp_54;
        end
        th_comp_54: begin
          th_comp <= th_comp_55;
        end
        th_comp_55: begin
          th_comp <= th_comp_56;
        end
        th_comp_56: begin
          th_comp <= th_comp_57;
        end
        th_comp_57: begin
          th_comp <= th_comp_58;
        end
        th_comp_58: begin
          th_comp <= th_comp_59;
        end
        th_comp_59: begin
          th_comp <= th_comp_60;
        end
        th_comp_60: begin
          th_comp <= th_comp_61;
        end
        th_comp_61: begin
          th_comp <= th_comp_62;
        end
        th_comp_62: begin
          th_comp <= th_comp_63;
        end
        th_comp_63: begin
          th_comp <= th_comp_64;
        end
        th_comp_64: begin
          th_comp <= th_comp_65;
        end
        th_comp_65: begin
          th_comp <= th_comp_66;
        end
        th_comp_66: begin
          th_comp <= th_comp_67;
        end
        th_comp_67: begin
          th_comp <= th_comp_68;
        end
        th_comp_68: begin
          th_comp <= th_comp_69;
        end
        th_comp_69: begin
          th_comp <= th_comp_70;
        end
        th_comp_70: begin
          th_comp <= th_comp_71;
        end
        th_comp_71: begin
          th_comp <= th_comp_72;
        end
        th_comp_72: begin
          th_comp <= th_comp_73;
        end
        th_comp_73: begin
          th_comp <= th_comp_74;
        end
        th_comp_74: begin
          th_comp <= th_comp_75;
        end
        th_comp_75: begin
          th_comp <= th_comp_76;
        end
        th_comp_76: begin
          th_comp <= th_comp_77;
        end
        th_comp_77: begin
          th_comp <= th_comp_78;
        end
        th_comp_78: begin
          th_comp <= th_comp_79;
        end
        th_comp_79: begin
          th_comp <= th_comp_80;
        end
        th_comp_80: begin
          _th_comp_end_time_6 <= counter;
          th_comp <= th_comp_81;
        end
        th_comp_81: begin
          $display("# para = %d, exec2_time = %d", 32, (_th_comp_end_time_6 - _th_comp_start_time_5));
          th_comp <= th_comp_82;
        end
        th_comp_82: begin
          _th_comp_end_time_6 <= counter;
          th_comp <= th_comp_83;
        end
        th_comp_83: begin
          $display("# para = %d, exec_time = %d", 32, (_th_comp_end_time_6 - _th_comp_start_time_5));
          th_comp <= th_comp_84;
        end
        th_comp_84: begin
          th_comp <= th_comp_85;
        end
        th_comp_85: begin
          if(_mystream_busy) begin
            th_comp <= th_comp_86;
          end 
        end
        th_comp_86: begin
          if(!_mystream_busy) begin
            th_comp <= th_comp_87;
          end 
        end
        th_comp_87: begin
          _th_comp_end_time_6 <= counter;
          th_comp <= th_comp_88;
        end
        th_comp_88: begin
          _th_comp_exec_time_7 <= _th_comp_end_time_6 - _th_comp_start_time_5;
          th_comp <= th_comp_89;
        end
        th_comp_89: begin
          $display("# para = %d, exec_time = %d", 32, _th_comp_exec_time_7);
          th_comp <= th_comp_90;
        end
        th_comp_90: begin
          _th_comp_offset_2 <= 512;
          th_comp <= th_comp_91;
        end
        th_comp_91: begin
          if(_myaxi_read_req_idle) begin
            th_comp <= th_comp_92;
          end 
        end
        th_comp_92: begin
          if(_myaxi_read_idle) begin
            th_comp <= th_comp_93;
          end 
        end
        th_comp_93: begin
          if(_myaxi_read_req_idle) begin
            th_comp <= th_comp_94;
          end 
        end
        th_comp_94: begin
          if(_myaxi_read_idle) begin
            th_comp <= th_comp_95;
          end 
        end
        th_comp_95: begin
          _th_comp_size_8 <= _th_comp_size_0;
          _th_comp_offset_9 <= _th_comp_offset_2;
          th_comp <= th_comp_96;
        end
        th_comp_96: begin
          _th_comp_sum_10 <= 0;
          th_comp <= th_comp_97;
        end
        th_comp_97: begin
          _th_comp_i_11 <= 0;
          th_comp <= th_comp_98;
        end
        th_comp_98: begin
          if(_th_comp_i_11 < _th_comp_size_8) begin
            th_comp <= th_comp_99;
          end else begin
            th_comp <= th_comp_106;
          end
        end
        th_comp_99: begin
          if(__tmp_1098_1) begin
            read_rdata_1099 <= ram_x_0_rdata;
          end 
          if(__tmp_1098_1) begin
            th_comp <= th_comp_100;
          end 
        end
        th_comp_100: begin
          _th_comp_a_12 <= read_rdata_1099;
          th_comp <= th_comp_101;
        end
        th_comp_101: begin
          if(__tmp_1101_1) begin
            read_rdata_1102 <= ram_y_0_rdata;
          end 
          if(__tmp_1101_1) begin
            th_comp <= th_comp_102;
          end 
        end
        th_comp_102: begin
          _th_comp_b_13 <= read_rdata_1102;
          th_comp <= th_comp_103;
        end
        th_comp_103: begin
          _th_comp_sum_10 <= _th_comp_a_12 + _th_comp_b_13;
          th_comp <= th_comp_104;
        end
        th_comp_104: begin
          th_comp <= th_comp_105;
        end
        th_comp_105: begin
          _th_comp_i_11 <= _th_comp_i_11 + 1;
          th_comp <= th_comp_98;
        end
        th_comp_106: begin
          if(_myaxi_write_req_idle) begin
            th_comp <= th_comp_107;
          end 
        end
        th_comp_107: begin
          if(_myaxi_write_idle && (outstanding_wcount_0 == 0)) begin
            th_comp <= th_comp_108;
          end 
        end
        th_comp_108: begin
          if(_myaxi_read_req_idle) begin
            th_comp <= th_comp_109;
          end 
        end
        th_comp_109: begin
          if(_myaxi_read_idle) begin
            th_comp <= th_comp_110;
          end 
        end
        th_comp_110: begin
          _th_comp_size_14 <= _th_comp_size_0;
          _th_comp_offset_stream_15 <= 0;
          _th_comp_offset_seq_16 <= _th_comp_offset_2;
          th_comp <= th_comp_111;
        end
        th_comp_111: begin
          _th_comp_all_ok_17 <= 1;
          th_comp <= th_comp_112;
        end
        th_comp_112: begin
          _th_comp_i_18 <= 0;
          th_comp <= th_comp_113;
        end
        th_comp_113: begin
          if(_th_comp_i_18 < _th_comp_size_14) begin
            th_comp <= th_comp_114;
          end else begin
            th_comp <= th_comp_121;
          end
        end
        th_comp_114: begin
          if(read_rtl_rvalid_1284) begin
            read_rdata_1285 <= read_rtl_rdata_1283;
          end 
          if(read_rtl_rvalid_1284) begin
            th_comp <= th_comp_115;
          end 
        end
        th_comp_115: begin
          _th_comp_st_19 <= read_rdata_1285;
          th_comp <= th_comp_116;
        end
        th_comp_116: begin
          if(read_rtl_rvalid_1353) begin
            read_rdata_1354 <= read_rtl_rdata_1352;
          end 
          if(read_rtl_rvalid_1353) begin
            th_comp <= th_comp_117;
          end 
        end
        th_comp_117: begin
          _th_comp_sq_20 <= read_rdata_1354;
          th_comp <= th_comp_118;
        end
        th_comp_118: begin
          if(_th_comp_st_19 !== _th_comp_sq_20) begin
            th_comp <= th_comp_119;
          end else begin
            th_comp <= th_comp_120;
          end
        end
        th_comp_119: begin
          _th_comp_all_ok_17 <= 0;
          th_comp <= th_comp_120;
        end
        th_comp_120: begin
          _th_comp_i_18 <= _th_comp_i_18 + 1;
          th_comp <= th_comp_113;
        end
        th_comp_121: begin
          if(_th_comp_all_ok_17) begin
            th_comp <= th_comp_122;
          end else begin
            th_comp <= th_comp_124;
          end
        end
        th_comp_122: begin
          $display("# verify: PASSED");
          th_comp <= th_comp_123;
        end
        th_comp_123: begin
          th_comp <= th_comp_125;
        end
        th_comp_124: begin
          $display("# verify: FAILED");
          th_comp <= th_comp_125;
        end
        th_comp_125: begin
          $finish;
          th_comp <= th_comp_126;
        end
      endcase
    end
  end

  localparam _myaxi_read_req_fsm_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      _myaxi_read_req_fsm <= _myaxi_read_req_fsm_init;
      _myaxi_read_cont <= 0;
    end else begin
      case(_myaxi_read_req_fsm)
        _myaxi_read_req_fsm_init: begin
          if((_myaxi_read_req_fsm == 0) && (_myaxi_read_start || _myaxi_read_cont) && !_myaxi_read_req_fifo_almost_full) begin
            _myaxi_read_req_fsm <= _myaxi_read_req_fsm_1;
          end 
        end
        _myaxi_read_req_fsm_1: begin
          if(myaxi_arready || !myaxi_arvalid) begin
            _myaxi_read_cont <= 1;
          end 
          if((myaxi_arready || !myaxi_arvalid) && (_myaxi_read_global_size == 0)) begin
            _myaxi_read_cont <= 0;
          end 
          if(myaxi_arready || !myaxi_arvalid) begin
            _myaxi_read_req_fsm <= _myaxi_read_req_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam _myaxi_read_data_narrow_fsm_1 = 1;
  localparam _myaxi_read_data_narrow_fsm_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _myaxi_read_data_narrow_fsm <= _myaxi_read_data_narrow_fsm_init;
      _myaxi_read_narrow_count_38 <= 0;
      _myaxi_read_narrow_wvalid_37 <= 0;
      _myaxi_read_narrow_wdata_36 <= 0;
      _myaxi_read_narrow_count_114 <= 0;
      _myaxi_read_narrow_wvalid_113 <= 0;
      _myaxi_read_narrow_wdata_112 <= 0;
      _myaxi_read_narrow_count_1148 <= 0;
      _myaxi_read_narrow_wvalid_1147 <= 0;
      _myaxi_read_narrow_wdata_1146 <= 0;
    end else begin
      case(_myaxi_read_data_narrow_fsm)
        _myaxi_read_data_narrow_fsm_init: begin
          if(_myaxi_read_data_idle && !_myaxi_read_req_fifo_empty && (_myaxi_read_op_sel_fifo == 1)) begin
            _myaxi_read_data_narrow_fsm <= _myaxi_read_data_narrow_fsm_1;
          end 
          if(_myaxi_read_data_idle && !_myaxi_read_req_fifo_empty && (_myaxi_read_op_sel_fifo == 2)) begin
            _myaxi_read_data_narrow_fsm <= _myaxi_read_data_narrow_fsm_1;
          end 
          if(_myaxi_read_data_idle && !_myaxi_read_req_fifo_empty && (_myaxi_read_op_sel_fifo == 5)) begin
            _myaxi_read_data_narrow_fsm <= _myaxi_read_data_narrow_fsm_1;
          end 
        end
        _myaxi_read_data_narrow_fsm_1: begin
          _myaxi_read_narrow_count_38 <= 0;
          _myaxi_read_narrow_wvalid_37 <= 0;
          _myaxi_read_narrow_count_114 <= 0;
          _myaxi_read_narrow_wvalid_113 <= 0;
          _myaxi_read_narrow_count_1148 <= 0;
          _myaxi_read_narrow_wvalid_1147 <= 0;
          _myaxi_read_data_narrow_fsm <= _myaxi_read_data_narrow_fsm_2;
          _myaxi_read_data_narrow_fsm <= _myaxi_read_data_narrow_fsm_2;
          _myaxi_read_data_narrow_fsm <= _myaxi_read_data_narrow_fsm_2;
        end
        _myaxi_read_data_narrow_fsm_2: begin
          if(_myaxi_read_op_sel_buf == 1) begin
            _myaxi_read_narrow_wvalid_37 <= 0;
          end 
          if((_myaxi_read_op_sel_buf == 1) && myaxi_rvalid && (_myaxi_read_narrow_count_38 < 31)) begin
            _myaxi_read_narrow_count_38 <= _myaxi_read_narrow_count_38 + 1;
            _myaxi_read_narrow_wdata_36 <= { myaxi_rdata, _myaxi_read_narrow_wdata_36[1023:32] };
            _myaxi_read_narrow_wvalid_37 <= 0;
          end 
          if((_myaxi_read_op_sel_buf == 1) && myaxi_rvalid && (_myaxi_read_narrow_count_38 == 31)) begin
            _myaxi_read_narrow_count_38 <= 0;
            _myaxi_read_narrow_wdata_36 <= { myaxi_rdata, _myaxi_read_narrow_wdata_36[1023:32] };
            _myaxi_read_narrow_wvalid_37 <= 1;
          end 
          if(_myaxi_read_op_sel_buf == 2) begin
            _myaxi_read_narrow_wvalid_113 <= 0;
          end 
          if((_myaxi_read_op_sel_buf == 2) && myaxi_rvalid && (_myaxi_read_narrow_count_114 < 31)) begin
            _myaxi_read_narrow_count_114 <= _myaxi_read_narrow_count_114 + 1;
            _myaxi_read_narrow_wdata_112 <= { myaxi_rdata, _myaxi_read_narrow_wdata_112[1023:32] };
            _myaxi_read_narrow_wvalid_113 <= 0;
          end 
          if((_myaxi_read_op_sel_buf == 2) && myaxi_rvalid && (_myaxi_read_narrow_count_114 == 31)) begin
            _myaxi_read_narrow_count_114 <= 0;
            _myaxi_read_narrow_wdata_112 <= { myaxi_rdata, _myaxi_read_narrow_wdata_112[1023:32] };
            _myaxi_read_narrow_wvalid_113 <= 1;
          end 
          if(_myaxi_read_op_sel_buf == 5) begin
            _myaxi_read_narrow_wvalid_1147 <= 0;
          end 
          if((_myaxi_read_op_sel_buf == 5) && myaxi_rvalid && (_myaxi_read_narrow_count_1148 < 31)) begin
            _myaxi_read_narrow_count_1148 <= _myaxi_read_narrow_count_1148 + 1;
            _myaxi_read_narrow_wdata_1146 <= { myaxi_rdata, _myaxi_read_narrow_wdata_1146[1023:32] };
            _myaxi_read_narrow_wvalid_1147 <= 0;
          end 
          if((_myaxi_read_op_sel_buf == 5) && myaxi_rvalid && (_myaxi_read_narrow_count_1148 == 31)) begin
            _myaxi_read_narrow_count_1148 <= 0;
            _myaxi_read_narrow_wdata_1146 <= { myaxi_rdata, _myaxi_read_narrow_wdata_1146[1023:32] };
            _myaxi_read_narrow_wvalid_1147 <= 1;
          end 
          if((_myaxi_read_op_sel_buf == 1) && myaxi_rvalid && (_myaxi_read_local_size_buf <= 1) && (_myaxi_read_narrow_count_38 == 31)) begin
            _myaxi_read_data_narrow_fsm <= _myaxi_read_data_narrow_fsm_init;
          end 
          if((_myaxi_read_op_sel_buf == 2) && myaxi_rvalid && (_myaxi_read_local_size_buf <= 1) && (_myaxi_read_narrow_count_114 == 31)) begin
            _myaxi_read_data_narrow_fsm <= _myaxi_read_data_narrow_fsm_init;
          end 
          if((_myaxi_read_op_sel_buf == 5) && myaxi_rvalid && (_myaxi_read_local_size_buf <= 1) && (_myaxi_read_narrow_count_1148 == 31)) begin
            _myaxi_read_data_narrow_fsm <= _myaxi_read_data_narrow_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_0_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_0 <= write_burst_packed_fsm_0_init;
      write_burst_packed_addr_39 <= 0;
      write_burst_packed_stride_40 <= 0;
      write_burst_packed_length_41 <= 0;
      write_burst_packed_done_42 <= 0;
    end else begin
      case(write_burst_packed_fsm_0)
        write_burst_packed_fsm_0_init: begin
          write_burst_packed_addr_39 <= _myaxi_read_local_addr_buf;
          write_burst_packed_stride_40 <= _myaxi_read_local_stride_buf;
          write_burst_packed_length_41 <= _myaxi_read_local_size_buf;
          write_burst_packed_done_42 <= 0;
          if((_myaxi_read_data_narrow_fsm == 1) && (_myaxi_read_op_sel_buf == 1) && (_myaxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_0 <= write_burst_packed_fsm_0_1;
          end 
        end
        write_burst_packed_fsm_0_1: begin
          if(_myaxi_read_narrow_wvalid_37) begin
            write_burst_packed_addr_39 <= write_burst_packed_addr_39 + write_burst_packed_stride_40;
            write_burst_packed_length_41 <= write_burst_packed_length_41 - 1;
            write_burst_packed_done_42 <= 0;
          end 
          if(_myaxi_read_narrow_wvalid_37 && (write_burst_packed_length_41 <= 1)) begin
            write_burst_packed_done_42 <= 1;
          end 
          if(_myaxi_read_narrow_wvalid_37 && 0) begin
            write_burst_packed_done_42 <= 1;
          end 
          if(_myaxi_read_narrow_wvalid_37 && (write_burst_packed_length_41 <= 1)) begin
            write_burst_packed_fsm_0 <= write_burst_packed_fsm_0_init;
          end 
          if(_myaxi_read_narrow_wvalid_37 && 0) begin
            write_burst_packed_fsm_0 <= write_burst_packed_fsm_0_init;
          end 
          if(0) begin
            write_burst_packed_fsm_0 <= write_burst_packed_fsm_0_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_1_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_1 <= write_burst_packed_fsm_1_init;
      write_burst_packed_addr_115 <= 0;
      write_burst_packed_stride_116 <= 0;
      write_burst_packed_length_117 <= 0;
      write_burst_packed_done_118 <= 0;
    end else begin
      case(write_burst_packed_fsm_1)
        write_burst_packed_fsm_1_init: begin
          write_burst_packed_addr_115 <= _myaxi_read_local_addr_buf;
          write_burst_packed_stride_116 <= _myaxi_read_local_stride_buf;
          write_burst_packed_length_117 <= _myaxi_read_local_size_buf;
          write_burst_packed_done_118 <= 0;
          if((_myaxi_read_data_narrow_fsm == 1) && (_myaxi_read_op_sel_buf == 2) && (_myaxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_1 <= write_burst_packed_fsm_1_1;
          end 
        end
        write_burst_packed_fsm_1_1: begin
          if(_myaxi_read_narrow_wvalid_113) begin
            write_burst_packed_addr_115 <= write_burst_packed_addr_115 + write_burst_packed_stride_116;
            write_burst_packed_length_117 <= write_burst_packed_length_117 - 1;
            write_burst_packed_done_118 <= 0;
          end 
          if(_myaxi_read_narrow_wvalid_113 && (write_burst_packed_length_117 <= 1)) begin
            write_burst_packed_done_118 <= 1;
          end 
          if(_myaxi_read_narrow_wvalid_113 && 0) begin
            write_burst_packed_done_118 <= 1;
          end 
          if(_myaxi_read_narrow_wvalid_113 && (write_burst_packed_length_117 <= 1)) begin
            write_burst_packed_fsm_1 <= write_burst_packed_fsm_1_init;
          end 
          if(_myaxi_read_narrow_wvalid_113 && 0) begin
            write_burst_packed_fsm_1 <= write_burst_packed_fsm_1_init;
          end 
          if(0) begin
            write_burst_packed_fsm_1 <= write_burst_packed_fsm_1_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_a0_source_fsm_0_1 = 1;
  localparam _mystream_a0_source_fsm_0_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_a0_source_fsm_0 <= _mystream_a0_source_fsm_0_init;
    end else begin
      case(_mystream_a0_source_fsm_0)
        _mystream_a0_source_fsm_0_init: begin
          if(_mystream_source_start && _mystream_a0_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_a0_source_fsm_0 <= _mystream_a0_source_fsm_0_1;
          end 
        end
        _mystream_a0_source_fsm_0_1: begin
          if(_mystream_stream_oready) begin
            _mystream_a0_source_fsm_0 <= _mystream_a0_source_fsm_0_2;
          end 
        end
        _mystream_a0_source_fsm_0_2: begin
          if((_mystream_a0_source_count == 1) && _mystream_stream_oready) begin
            _mystream_a0_source_fsm_0 <= _mystream_a0_source_fsm_0_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_a0_source_fsm_0 <= _mystream_a0_source_fsm_0_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_a1_source_fsm_1_1 = 1;
  localparam _mystream_a1_source_fsm_1_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_a1_source_fsm_1 <= _mystream_a1_source_fsm_1_init;
    end else begin
      case(_mystream_a1_source_fsm_1)
        _mystream_a1_source_fsm_1_init: begin
          if(_mystream_source_start && _mystream_a1_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_a1_source_fsm_1 <= _mystream_a1_source_fsm_1_1;
          end 
        end
        _mystream_a1_source_fsm_1_1: begin
          if(_mystream_stream_oready) begin
            _mystream_a1_source_fsm_1 <= _mystream_a1_source_fsm_1_2;
          end 
        end
        _mystream_a1_source_fsm_1_2: begin
          if((_mystream_a1_source_count == 1) && _mystream_stream_oready) begin
            _mystream_a1_source_fsm_1 <= _mystream_a1_source_fsm_1_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_a1_source_fsm_1 <= _mystream_a1_source_fsm_1_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_a2_source_fsm_2_1 = 1;
  localparam _mystream_a2_source_fsm_2_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_a2_source_fsm_2 <= _mystream_a2_source_fsm_2_init;
    end else begin
      case(_mystream_a2_source_fsm_2)
        _mystream_a2_source_fsm_2_init: begin
          if(_mystream_source_start && _mystream_a2_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_a2_source_fsm_2 <= _mystream_a2_source_fsm_2_1;
          end 
        end
        _mystream_a2_source_fsm_2_1: begin
          if(_mystream_stream_oready) begin
            _mystream_a2_source_fsm_2 <= _mystream_a2_source_fsm_2_2;
          end 
        end
        _mystream_a2_source_fsm_2_2: begin
          if((_mystream_a2_source_count == 1) && _mystream_stream_oready) begin
            _mystream_a2_source_fsm_2 <= _mystream_a2_source_fsm_2_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_a2_source_fsm_2 <= _mystream_a2_source_fsm_2_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_a3_source_fsm_3_1 = 1;
  localparam _mystream_a3_source_fsm_3_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_a3_source_fsm_3 <= _mystream_a3_source_fsm_3_init;
    end else begin
      case(_mystream_a3_source_fsm_3)
        _mystream_a3_source_fsm_3_init: begin
          if(_mystream_source_start && _mystream_a3_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_a3_source_fsm_3 <= _mystream_a3_source_fsm_3_1;
          end 
        end
        _mystream_a3_source_fsm_3_1: begin
          if(_mystream_stream_oready) begin
            _mystream_a3_source_fsm_3 <= _mystream_a3_source_fsm_3_2;
          end 
        end
        _mystream_a3_source_fsm_3_2: begin
          if((_mystream_a3_source_count == 1) && _mystream_stream_oready) begin
            _mystream_a3_source_fsm_3 <= _mystream_a3_source_fsm_3_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_a3_source_fsm_3 <= _mystream_a3_source_fsm_3_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_a4_source_fsm_4_1 = 1;
  localparam _mystream_a4_source_fsm_4_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_a4_source_fsm_4 <= _mystream_a4_source_fsm_4_init;
    end else begin
      case(_mystream_a4_source_fsm_4)
        _mystream_a4_source_fsm_4_init: begin
          if(_mystream_source_start && _mystream_a4_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_a4_source_fsm_4 <= _mystream_a4_source_fsm_4_1;
          end 
        end
        _mystream_a4_source_fsm_4_1: begin
          if(_mystream_stream_oready) begin
            _mystream_a4_source_fsm_4 <= _mystream_a4_source_fsm_4_2;
          end 
        end
        _mystream_a4_source_fsm_4_2: begin
          if((_mystream_a4_source_count == 1) && _mystream_stream_oready) begin
            _mystream_a4_source_fsm_4 <= _mystream_a4_source_fsm_4_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_a4_source_fsm_4 <= _mystream_a4_source_fsm_4_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_a5_source_fsm_5_1 = 1;
  localparam _mystream_a5_source_fsm_5_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_a5_source_fsm_5 <= _mystream_a5_source_fsm_5_init;
    end else begin
      case(_mystream_a5_source_fsm_5)
        _mystream_a5_source_fsm_5_init: begin
          if(_mystream_source_start && _mystream_a5_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_a5_source_fsm_5 <= _mystream_a5_source_fsm_5_1;
          end 
        end
        _mystream_a5_source_fsm_5_1: begin
          if(_mystream_stream_oready) begin
            _mystream_a5_source_fsm_5 <= _mystream_a5_source_fsm_5_2;
          end 
        end
        _mystream_a5_source_fsm_5_2: begin
          if((_mystream_a5_source_count == 1) && _mystream_stream_oready) begin
            _mystream_a5_source_fsm_5 <= _mystream_a5_source_fsm_5_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_a5_source_fsm_5 <= _mystream_a5_source_fsm_5_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_a6_source_fsm_6_1 = 1;
  localparam _mystream_a6_source_fsm_6_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_a6_source_fsm_6 <= _mystream_a6_source_fsm_6_init;
    end else begin
      case(_mystream_a6_source_fsm_6)
        _mystream_a6_source_fsm_6_init: begin
          if(_mystream_source_start && _mystream_a6_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_a6_source_fsm_6 <= _mystream_a6_source_fsm_6_1;
          end 
        end
        _mystream_a6_source_fsm_6_1: begin
          if(_mystream_stream_oready) begin
            _mystream_a6_source_fsm_6 <= _mystream_a6_source_fsm_6_2;
          end 
        end
        _mystream_a6_source_fsm_6_2: begin
          if((_mystream_a6_source_count == 1) && _mystream_stream_oready) begin
            _mystream_a6_source_fsm_6 <= _mystream_a6_source_fsm_6_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_a6_source_fsm_6 <= _mystream_a6_source_fsm_6_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_a7_source_fsm_7_1 = 1;
  localparam _mystream_a7_source_fsm_7_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_a7_source_fsm_7 <= _mystream_a7_source_fsm_7_init;
    end else begin
      case(_mystream_a7_source_fsm_7)
        _mystream_a7_source_fsm_7_init: begin
          if(_mystream_source_start && _mystream_a7_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_a7_source_fsm_7 <= _mystream_a7_source_fsm_7_1;
          end 
        end
        _mystream_a7_source_fsm_7_1: begin
          if(_mystream_stream_oready) begin
            _mystream_a7_source_fsm_7 <= _mystream_a7_source_fsm_7_2;
          end 
        end
        _mystream_a7_source_fsm_7_2: begin
          if((_mystream_a7_source_count == 1) && _mystream_stream_oready) begin
            _mystream_a7_source_fsm_7 <= _mystream_a7_source_fsm_7_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_a7_source_fsm_7 <= _mystream_a7_source_fsm_7_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_a8_source_fsm_8_1 = 1;
  localparam _mystream_a8_source_fsm_8_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_a8_source_fsm_8 <= _mystream_a8_source_fsm_8_init;
    end else begin
      case(_mystream_a8_source_fsm_8)
        _mystream_a8_source_fsm_8_init: begin
          if(_mystream_source_start && _mystream_a8_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_a8_source_fsm_8 <= _mystream_a8_source_fsm_8_1;
          end 
        end
        _mystream_a8_source_fsm_8_1: begin
          if(_mystream_stream_oready) begin
            _mystream_a8_source_fsm_8 <= _mystream_a8_source_fsm_8_2;
          end 
        end
        _mystream_a8_source_fsm_8_2: begin
          if((_mystream_a8_source_count == 1) && _mystream_stream_oready) begin
            _mystream_a8_source_fsm_8 <= _mystream_a8_source_fsm_8_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_a8_source_fsm_8 <= _mystream_a8_source_fsm_8_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_a9_source_fsm_9_1 = 1;
  localparam _mystream_a9_source_fsm_9_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_a9_source_fsm_9 <= _mystream_a9_source_fsm_9_init;
    end else begin
      case(_mystream_a9_source_fsm_9)
        _mystream_a9_source_fsm_9_init: begin
          if(_mystream_source_start && _mystream_a9_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_a9_source_fsm_9 <= _mystream_a9_source_fsm_9_1;
          end 
        end
        _mystream_a9_source_fsm_9_1: begin
          if(_mystream_stream_oready) begin
            _mystream_a9_source_fsm_9 <= _mystream_a9_source_fsm_9_2;
          end 
        end
        _mystream_a9_source_fsm_9_2: begin
          if((_mystream_a9_source_count == 1) && _mystream_stream_oready) begin
            _mystream_a9_source_fsm_9 <= _mystream_a9_source_fsm_9_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_a9_source_fsm_9 <= _mystream_a9_source_fsm_9_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_a10_source_fsm_10_1 = 1;
  localparam _mystream_a10_source_fsm_10_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_a10_source_fsm_10 <= _mystream_a10_source_fsm_10_init;
    end else begin
      case(_mystream_a10_source_fsm_10)
        _mystream_a10_source_fsm_10_init: begin
          if(_mystream_source_start && _mystream_a10_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_a10_source_fsm_10 <= _mystream_a10_source_fsm_10_1;
          end 
        end
        _mystream_a10_source_fsm_10_1: begin
          if(_mystream_stream_oready) begin
            _mystream_a10_source_fsm_10 <= _mystream_a10_source_fsm_10_2;
          end 
        end
        _mystream_a10_source_fsm_10_2: begin
          if((_mystream_a10_source_count == 1) && _mystream_stream_oready) begin
            _mystream_a10_source_fsm_10 <= _mystream_a10_source_fsm_10_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_a10_source_fsm_10 <= _mystream_a10_source_fsm_10_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_a11_source_fsm_11_1 = 1;
  localparam _mystream_a11_source_fsm_11_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_a11_source_fsm_11 <= _mystream_a11_source_fsm_11_init;
    end else begin
      case(_mystream_a11_source_fsm_11)
        _mystream_a11_source_fsm_11_init: begin
          if(_mystream_source_start && _mystream_a11_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_a11_source_fsm_11 <= _mystream_a11_source_fsm_11_1;
          end 
        end
        _mystream_a11_source_fsm_11_1: begin
          if(_mystream_stream_oready) begin
            _mystream_a11_source_fsm_11 <= _mystream_a11_source_fsm_11_2;
          end 
        end
        _mystream_a11_source_fsm_11_2: begin
          if((_mystream_a11_source_count == 1) && _mystream_stream_oready) begin
            _mystream_a11_source_fsm_11 <= _mystream_a11_source_fsm_11_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_a11_source_fsm_11 <= _mystream_a11_source_fsm_11_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_a12_source_fsm_12_1 = 1;
  localparam _mystream_a12_source_fsm_12_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_a12_source_fsm_12 <= _mystream_a12_source_fsm_12_init;
    end else begin
      case(_mystream_a12_source_fsm_12)
        _mystream_a12_source_fsm_12_init: begin
          if(_mystream_source_start && _mystream_a12_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_a12_source_fsm_12 <= _mystream_a12_source_fsm_12_1;
          end 
        end
        _mystream_a12_source_fsm_12_1: begin
          if(_mystream_stream_oready) begin
            _mystream_a12_source_fsm_12 <= _mystream_a12_source_fsm_12_2;
          end 
        end
        _mystream_a12_source_fsm_12_2: begin
          if((_mystream_a12_source_count == 1) && _mystream_stream_oready) begin
            _mystream_a12_source_fsm_12 <= _mystream_a12_source_fsm_12_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_a12_source_fsm_12 <= _mystream_a12_source_fsm_12_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_a13_source_fsm_13_1 = 1;
  localparam _mystream_a13_source_fsm_13_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_a13_source_fsm_13 <= _mystream_a13_source_fsm_13_init;
    end else begin
      case(_mystream_a13_source_fsm_13)
        _mystream_a13_source_fsm_13_init: begin
          if(_mystream_source_start && _mystream_a13_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_a13_source_fsm_13 <= _mystream_a13_source_fsm_13_1;
          end 
        end
        _mystream_a13_source_fsm_13_1: begin
          if(_mystream_stream_oready) begin
            _mystream_a13_source_fsm_13 <= _mystream_a13_source_fsm_13_2;
          end 
        end
        _mystream_a13_source_fsm_13_2: begin
          if((_mystream_a13_source_count == 1) && _mystream_stream_oready) begin
            _mystream_a13_source_fsm_13 <= _mystream_a13_source_fsm_13_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_a13_source_fsm_13 <= _mystream_a13_source_fsm_13_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_a14_source_fsm_14_1 = 1;
  localparam _mystream_a14_source_fsm_14_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_a14_source_fsm_14 <= _mystream_a14_source_fsm_14_init;
    end else begin
      case(_mystream_a14_source_fsm_14)
        _mystream_a14_source_fsm_14_init: begin
          if(_mystream_source_start && _mystream_a14_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_a14_source_fsm_14 <= _mystream_a14_source_fsm_14_1;
          end 
        end
        _mystream_a14_source_fsm_14_1: begin
          if(_mystream_stream_oready) begin
            _mystream_a14_source_fsm_14 <= _mystream_a14_source_fsm_14_2;
          end 
        end
        _mystream_a14_source_fsm_14_2: begin
          if((_mystream_a14_source_count == 1) && _mystream_stream_oready) begin
            _mystream_a14_source_fsm_14 <= _mystream_a14_source_fsm_14_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_a14_source_fsm_14 <= _mystream_a14_source_fsm_14_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_a15_source_fsm_15_1 = 1;
  localparam _mystream_a15_source_fsm_15_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_a15_source_fsm_15 <= _mystream_a15_source_fsm_15_init;
    end else begin
      case(_mystream_a15_source_fsm_15)
        _mystream_a15_source_fsm_15_init: begin
          if(_mystream_source_start && _mystream_a15_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_a15_source_fsm_15 <= _mystream_a15_source_fsm_15_1;
          end 
        end
        _mystream_a15_source_fsm_15_1: begin
          if(_mystream_stream_oready) begin
            _mystream_a15_source_fsm_15 <= _mystream_a15_source_fsm_15_2;
          end 
        end
        _mystream_a15_source_fsm_15_2: begin
          if((_mystream_a15_source_count == 1) && _mystream_stream_oready) begin
            _mystream_a15_source_fsm_15 <= _mystream_a15_source_fsm_15_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_a15_source_fsm_15 <= _mystream_a15_source_fsm_15_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_a16_source_fsm_16_1 = 1;
  localparam _mystream_a16_source_fsm_16_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_a16_source_fsm_16 <= _mystream_a16_source_fsm_16_init;
    end else begin
      case(_mystream_a16_source_fsm_16)
        _mystream_a16_source_fsm_16_init: begin
          if(_mystream_source_start && _mystream_a16_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_a16_source_fsm_16 <= _mystream_a16_source_fsm_16_1;
          end 
        end
        _mystream_a16_source_fsm_16_1: begin
          if(_mystream_stream_oready) begin
            _mystream_a16_source_fsm_16 <= _mystream_a16_source_fsm_16_2;
          end 
        end
        _mystream_a16_source_fsm_16_2: begin
          if((_mystream_a16_source_count == 1) && _mystream_stream_oready) begin
            _mystream_a16_source_fsm_16 <= _mystream_a16_source_fsm_16_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_a16_source_fsm_16 <= _mystream_a16_source_fsm_16_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_a17_source_fsm_17_1 = 1;
  localparam _mystream_a17_source_fsm_17_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_a17_source_fsm_17 <= _mystream_a17_source_fsm_17_init;
    end else begin
      case(_mystream_a17_source_fsm_17)
        _mystream_a17_source_fsm_17_init: begin
          if(_mystream_source_start && _mystream_a17_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_a17_source_fsm_17 <= _mystream_a17_source_fsm_17_1;
          end 
        end
        _mystream_a17_source_fsm_17_1: begin
          if(_mystream_stream_oready) begin
            _mystream_a17_source_fsm_17 <= _mystream_a17_source_fsm_17_2;
          end 
        end
        _mystream_a17_source_fsm_17_2: begin
          if((_mystream_a17_source_count == 1) && _mystream_stream_oready) begin
            _mystream_a17_source_fsm_17 <= _mystream_a17_source_fsm_17_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_a17_source_fsm_17 <= _mystream_a17_source_fsm_17_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_a18_source_fsm_18_1 = 1;
  localparam _mystream_a18_source_fsm_18_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_a18_source_fsm_18 <= _mystream_a18_source_fsm_18_init;
    end else begin
      case(_mystream_a18_source_fsm_18)
        _mystream_a18_source_fsm_18_init: begin
          if(_mystream_source_start && _mystream_a18_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_a18_source_fsm_18 <= _mystream_a18_source_fsm_18_1;
          end 
        end
        _mystream_a18_source_fsm_18_1: begin
          if(_mystream_stream_oready) begin
            _mystream_a18_source_fsm_18 <= _mystream_a18_source_fsm_18_2;
          end 
        end
        _mystream_a18_source_fsm_18_2: begin
          if((_mystream_a18_source_count == 1) && _mystream_stream_oready) begin
            _mystream_a18_source_fsm_18 <= _mystream_a18_source_fsm_18_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_a18_source_fsm_18 <= _mystream_a18_source_fsm_18_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_a19_source_fsm_19_1 = 1;
  localparam _mystream_a19_source_fsm_19_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_a19_source_fsm_19 <= _mystream_a19_source_fsm_19_init;
    end else begin
      case(_mystream_a19_source_fsm_19)
        _mystream_a19_source_fsm_19_init: begin
          if(_mystream_source_start && _mystream_a19_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_a19_source_fsm_19 <= _mystream_a19_source_fsm_19_1;
          end 
        end
        _mystream_a19_source_fsm_19_1: begin
          if(_mystream_stream_oready) begin
            _mystream_a19_source_fsm_19 <= _mystream_a19_source_fsm_19_2;
          end 
        end
        _mystream_a19_source_fsm_19_2: begin
          if((_mystream_a19_source_count == 1) && _mystream_stream_oready) begin
            _mystream_a19_source_fsm_19 <= _mystream_a19_source_fsm_19_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_a19_source_fsm_19 <= _mystream_a19_source_fsm_19_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_a20_source_fsm_20_1 = 1;
  localparam _mystream_a20_source_fsm_20_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_a20_source_fsm_20 <= _mystream_a20_source_fsm_20_init;
    end else begin
      case(_mystream_a20_source_fsm_20)
        _mystream_a20_source_fsm_20_init: begin
          if(_mystream_source_start && _mystream_a20_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_a20_source_fsm_20 <= _mystream_a20_source_fsm_20_1;
          end 
        end
        _mystream_a20_source_fsm_20_1: begin
          if(_mystream_stream_oready) begin
            _mystream_a20_source_fsm_20 <= _mystream_a20_source_fsm_20_2;
          end 
        end
        _mystream_a20_source_fsm_20_2: begin
          if((_mystream_a20_source_count == 1) && _mystream_stream_oready) begin
            _mystream_a20_source_fsm_20 <= _mystream_a20_source_fsm_20_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_a20_source_fsm_20 <= _mystream_a20_source_fsm_20_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_a21_source_fsm_21_1 = 1;
  localparam _mystream_a21_source_fsm_21_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_a21_source_fsm_21 <= _mystream_a21_source_fsm_21_init;
    end else begin
      case(_mystream_a21_source_fsm_21)
        _mystream_a21_source_fsm_21_init: begin
          if(_mystream_source_start && _mystream_a21_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_a21_source_fsm_21 <= _mystream_a21_source_fsm_21_1;
          end 
        end
        _mystream_a21_source_fsm_21_1: begin
          if(_mystream_stream_oready) begin
            _mystream_a21_source_fsm_21 <= _mystream_a21_source_fsm_21_2;
          end 
        end
        _mystream_a21_source_fsm_21_2: begin
          if((_mystream_a21_source_count == 1) && _mystream_stream_oready) begin
            _mystream_a21_source_fsm_21 <= _mystream_a21_source_fsm_21_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_a21_source_fsm_21 <= _mystream_a21_source_fsm_21_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_a22_source_fsm_22_1 = 1;
  localparam _mystream_a22_source_fsm_22_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_a22_source_fsm_22 <= _mystream_a22_source_fsm_22_init;
    end else begin
      case(_mystream_a22_source_fsm_22)
        _mystream_a22_source_fsm_22_init: begin
          if(_mystream_source_start && _mystream_a22_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_a22_source_fsm_22 <= _mystream_a22_source_fsm_22_1;
          end 
        end
        _mystream_a22_source_fsm_22_1: begin
          if(_mystream_stream_oready) begin
            _mystream_a22_source_fsm_22 <= _mystream_a22_source_fsm_22_2;
          end 
        end
        _mystream_a22_source_fsm_22_2: begin
          if((_mystream_a22_source_count == 1) && _mystream_stream_oready) begin
            _mystream_a22_source_fsm_22 <= _mystream_a22_source_fsm_22_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_a22_source_fsm_22 <= _mystream_a22_source_fsm_22_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_a23_source_fsm_23_1 = 1;
  localparam _mystream_a23_source_fsm_23_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_a23_source_fsm_23 <= _mystream_a23_source_fsm_23_init;
    end else begin
      case(_mystream_a23_source_fsm_23)
        _mystream_a23_source_fsm_23_init: begin
          if(_mystream_source_start && _mystream_a23_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_a23_source_fsm_23 <= _mystream_a23_source_fsm_23_1;
          end 
        end
        _mystream_a23_source_fsm_23_1: begin
          if(_mystream_stream_oready) begin
            _mystream_a23_source_fsm_23 <= _mystream_a23_source_fsm_23_2;
          end 
        end
        _mystream_a23_source_fsm_23_2: begin
          if((_mystream_a23_source_count == 1) && _mystream_stream_oready) begin
            _mystream_a23_source_fsm_23 <= _mystream_a23_source_fsm_23_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_a23_source_fsm_23 <= _mystream_a23_source_fsm_23_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_a24_source_fsm_24_1 = 1;
  localparam _mystream_a24_source_fsm_24_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_a24_source_fsm_24 <= _mystream_a24_source_fsm_24_init;
    end else begin
      case(_mystream_a24_source_fsm_24)
        _mystream_a24_source_fsm_24_init: begin
          if(_mystream_source_start && _mystream_a24_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_a24_source_fsm_24 <= _mystream_a24_source_fsm_24_1;
          end 
        end
        _mystream_a24_source_fsm_24_1: begin
          if(_mystream_stream_oready) begin
            _mystream_a24_source_fsm_24 <= _mystream_a24_source_fsm_24_2;
          end 
        end
        _mystream_a24_source_fsm_24_2: begin
          if((_mystream_a24_source_count == 1) && _mystream_stream_oready) begin
            _mystream_a24_source_fsm_24 <= _mystream_a24_source_fsm_24_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_a24_source_fsm_24 <= _mystream_a24_source_fsm_24_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_a25_source_fsm_25_1 = 1;
  localparam _mystream_a25_source_fsm_25_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_a25_source_fsm_25 <= _mystream_a25_source_fsm_25_init;
    end else begin
      case(_mystream_a25_source_fsm_25)
        _mystream_a25_source_fsm_25_init: begin
          if(_mystream_source_start && _mystream_a25_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_a25_source_fsm_25 <= _mystream_a25_source_fsm_25_1;
          end 
        end
        _mystream_a25_source_fsm_25_1: begin
          if(_mystream_stream_oready) begin
            _mystream_a25_source_fsm_25 <= _mystream_a25_source_fsm_25_2;
          end 
        end
        _mystream_a25_source_fsm_25_2: begin
          if((_mystream_a25_source_count == 1) && _mystream_stream_oready) begin
            _mystream_a25_source_fsm_25 <= _mystream_a25_source_fsm_25_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_a25_source_fsm_25 <= _mystream_a25_source_fsm_25_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_a26_source_fsm_26_1 = 1;
  localparam _mystream_a26_source_fsm_26_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_a26_source_fsm_26 <= _mystream_a26_source_fsm_26_init;
    end else begin
      case(_mystream_a26_source_fsm_26)
        _mystream_a26_source_fsm_26_init: begin
          if(_mystream_source_start && _mystream_a26_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_a26_source_fsm_26 <= _mystream_a26_source_fsm_26_1;
          end 
        end
        _mystream_a26_source_fsm_26_1: begin
          if(_mystream_stream_oready) begin
            _mystream_a26_source_fsm_26 <= _mystream_a26_source_fsm_26_2;
          end 
        end
        _mystream_a26_source_fsm_26_2: begin
          if((_mystream_a26_source_count == 1) && _mystream_stream_oready) begin
            _mystream_a26_source_fsm_26 <= _mystream_a26_source_fsm_26_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_a26_source_fsm_26 <= _mystream_a26_source_fsm_26_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_a27_source_fsm_27_1 = 1;
  localparam _mystream_a27_source_fsm_27_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_a27_source_fsm_27 <= _mystream_a27_source_fsm_27_init;
    end else begin
      case(_mystream_a27_source_fsm_27)
        _mystream_a27_source_fsm_27_init: begin
          if(_mystream_source_start && _mystream_a27_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_a27_source_fsm_27 <= _mystream_a27_source_fsm_27_1;
          end 
        end
        _mystream_a27_source_fsm_27_1: begin
          if(_mystream_stream_oready) begin
            _mystream_a27_source_fsm_27 <= _mystream_a27_source_fsm_27_2;
          end 
        end
        _mystream_a27_source_fsm_27_2: begin
          if((_mystream_a27_source_count == 1) && _mystream_stream_oready) begin
            _mystream_a27_source_fsm_27 <= _mystream_a27_source_fsm_27_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_a27_source_fsm_27 <= _mystream_a27_source_fsm_27_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_a28_source_fsm_28_1 = 1;
  localparam _mystream_a28_source_fsm_28_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_a28_source_fsm_28 <= _mystream_a28_source_fsm_28_init;
    end else begin
      case(_mystream_a28_source_fsm_28)
        _mystream_a28_source_fsm_28_init: begin
          if(_mystream_source_start && _mystream_a28_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_a28_source_fsm_28 <= _mystream_a28_source_fsm_28_1;
          end 
        end
        _mystream_a28_source_fsm_28_1: begin
          if(_mystream_stream_oready) begin
            _mystream_a28_source_fsm_28 <= _mystream_a28_source_fsm_28_2;
          end 
        end
        _mystream_a28_source_fsm_28_2: begin
          if((_mystream_a28_source_count == 1) && _mystream_stream_oready) begin
            _mystream_a28_source_fsm_28 <= _mystream_a28_source_fsm_28_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_a28_source_fsm_28 <= _mystream_a28_source_fsm_28_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_a29_source_fsm_29_1 = 1;
  localparam _mystream_a29_source_fsm_29_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_a29_source_fsm_29 <= _mystream_a29_source_fsm_29_init;
    end else begin
      case(_mystream_a29_source_fsm_29)
        _mystream_a29_source_fsm_29_init: begin
          if(_mystream_source_start && _mystream_a29_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_a29_source_fsm_29 <= _mystream_a29_source_fsm_29_1;
          end 
        end
        _mystream_a29_source_fsm_29_1: begin
          if(_mystream_stream_oready) begin
            _mystream_a29_source_fsm_29 <= _mystream_a29_source_fsm_29_2;
          end 
        end
        _mystream_a29_source_fsm_29_2: begin
          if((_mystream_a29_source_count == 1) && _mystream_stream_oready) begin
            _mystream_a29_source_fsm_29 <= _mystream_a29_source_fsm_29_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_a29_source_fsm_29 <= _mystream_a29_source_fsm_29_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_a30_source_fsm_30_1 = 1;
  localparam _mystream_a30_source_fsm_30_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_a30_source_fsm_30 <= _mystream_a30_source_fsm_30_init;
    end else begin
      case(_mystream_a30_source_fsm_30)
        _mystream_a30_source_fsm_30_init: begin
          if(_mystream_source_start && _mystream_a30_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_a30_source_fsm_30 <= _mystream_a30_source_fsm_30_1;
          end 
        end
        _mystream_a30_source_fsm_30_1: begin
          if(_mystream_stream_oready) begin
            _mystream_a30_source_fsm_30 <= _mystream_a30_source_fsm_30_2;
          end 
        end
        _mystream_a30_source_fsm_30_2: begin
          if((_mystream_a30_source_count == 1) && _mystream_stream_oready) begin
            _mystream_a30_source_fsm_30 <= _mystream_a30_source_fsm_30_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_a30_source_fsm_30 <= _mystream_a30_source_fsm_30_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_a31_source_fsm_31_1 = 1;
  localparam _mystream_a31_source_fsm_31_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_a31_source_fsm_31 <= _mystream_a31_source_fsm_31_init;
    end else begin
      case(_mystream_a31_source_fsm_31)
        _mystream_a31_source_fsm_31_init: begin
          if(_mystream_source_start && _mystream_a31_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_a31_source_fsm_31 <= _mystream_a31_source_fsm_31_1;
          end 
        end
        _mystream_a31_source_fsm_31_1: begin
          if(_mystream_stream_oready) begin
            _mystream_a31_source_fsm_31 <= _mystream_a31_source_fsm_31_2;
          end 
        end
        _mystream_a31_source_fsm_31_2: begin
          if((_mystream_a31_source_count == 1) && _mystream_stream_oready) begin
            _mystream_a31_source_fsm_31 <= _mystream_a31_source_fsm_31_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_a31_source_fsm_31 <= _mystream_a31_source_fsm_31_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_b0_source_fsm_32_1 = 1;
  localparam _mystream_b0_source_fsm_32_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_b0_source_fsm_32 <= _mystream_b0_source_fsm_32_init;
    end else begin
      case(_mystream_b0_source_fsm_32)
        _mystream_b0_source_fsm_32_init: begin
          if(_mystream_source_start && _mystream_b0_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_b0_source_fsm_32 <= _mystream_b0_source_fsm_32_1;
          end 
        end
        _mystream_b0_source_fsm_32_1: begin
          if(_mystream_stream_oready) begin
            _mystream_b0_source_fsm_32 <= _mystream_b0_source_fsm_32_2;
          end 
        end
        _mystream_b0_source_fsm_32_2: begin
          if((_mystream_b0_source_count == 1) && _mystream_stream_oready) begin
            _mystream_b0_source_fsm_32 <= _mystream_b0_source_fsm_32_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_b0_source_fsm_32 <= _mystream_b0_source_fsm_32_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_b1_source_fsm_33_1 = 1;
  localparam _mystream_b1_source_fsm_33_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_b1_source_fsm_33 <= _mystream_b1_source_fsm_33_init;
    end else begin
      case(_mystream_b1_source_fsm_33)
        _mystream_b1_source_fsm_33_init: begin
          if(_mystream_source_start && _mystream_b1_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_b1_source_fsm_33 <= _mystream_b1_source_fsm_33_1;
          end 
        end
        _mystream_b1_source_fsm_33_1: begin
          if(_mystream_stream_oready) begin
            _mystream_b1_source_fsm_33 <= _mystream_b1_source_fsm_33_2;
          end 
        end
        _mystream_b1_source_fsm_33_2: begin
          if((_mystream_b1_source_count == 1) && _mystream_stream_oready) begin
            _mystream_b1_source_fsm_33 <= _mystream_b1_source_fsm_33_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_b1_source_fsm_33 <= _mystream_b1_source_fsm_33_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_b2_source_fsm_34_1 = 1;
  localparam _mystream_b2_source_fsm_34_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_b2_source_fsm_34 <= _mystream_b2_source_fsm_34_init;
    end else begin
      case(_mystream_b2_source_fsm_34)
        _mystream_b2_source_fsm_34_init: begin
          if(_mystream_source_start && _mystream_b2_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_b2_source_fsm_34 <= _mystream_b2_source_fsm_34_1;
          end 
        end
        _mystream_b2_source_fsm_34_1: begin
          if(_mystream_stream_oready) begin
            _mystream_b2_source_fsm_34 <= _mystream_b2_source_fsm_34_2;
          end 
        end
        _mystream_b2_source_fsm_34_2: begin
          if((_mystream_b2_source_count == 1) && _mystream_stream_oready) begin
            _mystream_b2_source_fsm_34 <= _mystream_b2_source_fsm_34_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_b2_source_fsm_34 <= _mystream_b2_source_fsm_34_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_b3_source_fsm_35_1 = 1;
  localparam _mystream_b3_source_fsm_35_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_b3_source_fsm_35 <= _mystream_b3_source_fsm_35_init;
    end else begin
      case(_mystream_b3_source_fsm_35)
        _mystream_b3_source_fsm_35_init: begin
          if(_mystream_source_start && _mystream_b3_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_b3_source_fsm_35 <= _mystream_b3_source_fsm_35_1;
          end 
        end
        _mystream_b3_source_fsm_35_1: begin
          if(_mystream_stream_oready) begin
            _mystream_b3_source_fsm_35 <= _mystream_b3_source_fsm_35_2;
          end 
        end
        _mystream_b3_source_fsm_35_2: begin
          if((_mystream_b3_source_count == 1) && _mystream_stream_oready) begin
            _mystream_b3_source_fsm_35 <= _mystream_b3_source_fsm_35_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_b3_source_fsm_35 <= _mystream_b3_source_fsm_35_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_b4_source_fsm_36_1 = 1;
  localparam _mystream_b4_source_fsm_36_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_b4_source_fsm_36 <= _mystream_b4_source_fsm_36_init;
    end else begin
      case(_mystream_b4_source_fsm_36)
        _mystream_b4_source_fsm_36_init: begin
          if(_mystream_source_start && _mystream_b4_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_b4_source_fsm_36 <= _mystream_b4_source_fsm_36_1;
          end 
        end
        _mystream_b4_source_fsm_36_1: begin
          if(_mystream_stream_oready) begin
            _mystream_b4_source_fsm_36 <= _mystream_b4_source_fsm_36_2;
          end 
        end
        _mystream_b4_source_fsm_36_2: begin
          if((_mystream_b4_source_count == 1) && _mystream_stream_oready) begin
            _mystream_b4_source_fsm_36 <= _mystream_b4_source_fsm_36_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_b4_source_fsm_36 <= _mystream_b4_source_fsm_36_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_b5_source_fsm_37_1 = 1;
  localparam _mystream_b5_source_fsm_37_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_b5_source_fsm_37 <= _mystream_b5_source_fsm_37_init;
    end else begin
      case(_mystream_b5_source_fsm_37)
        _mystream_b5_source_fsm_37_init: begin
          if(_mystream_source_start && _mystream_b5_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_b5_source_fsm_37 <= _mystream_b5_source_fsm_37_1;
          end 
        end
        _mystream_b5_source_fsm_37_1: begin
          if(_mystream_stream_oready) begin
            _mystream_b5_source_fsm_37 <= _mystream_b5_source_fsm_37_2;
          end 
        end
        _mystream_b5_source_fsm_37_2: begin
          if((_mystream_b5_source_count == 1) && _mystream_stream_oready) begin
            _mystream_b5_source_fsm_37 <= _mystream_b5_source_fsm_37_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_b5_source_fsm_37 <= _mystream_b5_source_fsm_37_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_b6_source_fsm_38_1 = 1;
  localparam _mystream_b6_source_fsm_38_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_b6_source_fsm_38 <= _mystream_b6_source_fsm_38_init;
    end else begin
      case(_mystream_b6_source_fsm_38)
        _mystream_b6_source_fsm_38_init: begin
          if(_mystream_source_start && _mystream_b6_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_b6_source_fsm_38 <= _mystream_b6_source_fsm_38_1;
          end 
        end
        _mystream_b6_source_fsm_38_1: begin
          if(_mystream_stream_oready) begin
            _mystream_b6_source_fsm_38 <= _mystream_b6_source_fsm_38_2;
          end 
        end
        _mystream_b6_source_fsm_38_2: begin
          if((_mystream_b6_source_count == 1) && _mystream_stream_oready) begin
            _mystream_b6_source_fsm_38 <= _mystream_b6_source_fsm_38_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_b6_source_fsm_38 <= _mystream_b6_source_fsm_38_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_b7_source_fsm_39_1 = 1;
  localparam _mystream_b7_source_fsm_39_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_b7_source_fsm_39 <= _mystream_b7_source_fsm_39_init;
    end else begin
      case(_mystream_b7_source_fsm_39)
        _mystream_b7_source_fsm_39_init: begin
          if(_mystream_source_start && _mystream_b7_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_b7_source_fsm_39 <= _mystream_b7_source_fsm_39_1;
          end 
        end
        _mystream_b7_source_fsm_39_1: begin
          if(_mystream_stream_oready) begin
            _mystream_b7_source_fsm_39 <= _mystream_b7_source_fsm_39_2;
          end 
        end
        _mystream_b7_source_fsm_39_2: begin
          if((_mystream_b7_source_count == 1) && _mystream_stream_oready) begin
            _mystream_b7_source_fsm_39 <= _mystream_b7_source_fsm_39_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_b7_source_fsm_39 <= _mystream_b7_source_fsm_39_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_b8_source_fsm_40_1 = 1;
  localparam _mystream_b8_source_fsm_40_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_b8_source_fsm_40 <= _mystream_b8_source_fsm_40_init;
    end else begin
      case(_mystream_b8_source_fsm_40)
        _mystream_b8_source_fsm_40_init: begin
          if(_mystream_source_start && _mystream_b8_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_b8_source_fsm_40 <= _mystream_b8_source_fsm_40_1;
          end 
        end
        _mystream_b8_source_fsm_40_1: begin
          if(_mystream_stream_oready) begin
            _mystream_b8_source_fsm_40 <= _mystream_b8_source_fsm_40_2;
          end 
        end
        _mystream_b8_source_fsm_40_2: begin
          if((_mystream_b8_source_count == 1) && _mystream_stream_oready) begin
            _mystream_b8_source_fsm_40 <= _mystream_b8_source_fsm_40_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_b8_source_fsm_40 <= _mystream_b8_source_fsm_40_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_b9_source_fsm_41_1 = 1;
  localparam _mystream_b9_source_fsm_41_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_b9_source_fsm_41 <= _mystream_b9_source_fsm_41_init;
    end else begin
      case(_mystream_b9_source_fsm_41)
        _mystream_b9_source_fsm_41_init: begin
          if(_mystream_source_start && _mystream_b9_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_b9_source_fsm_41 <= _mystream_b9_source_fsm_41_1;
          end 
        end
        _mystream_b9_source_fsm_41_1: begin
          if(_mystream_stream_oready) begin
            _mystream_b9_source_fsm_41 <= _mystream_b9_source_fsm_41_2;
          end 
        end
        _mystream_b9_source_fsm_41_2: begin
          if((_mystream_b9_source_count == 1) && _mystream_stream_oready) begin
            _mystream_b9_source_fsm_41 <= _mystream_b9_source_fsm_41_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_b9_source_fsm_41 <= _mystream_b9_source_fsm_41_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_b10_source_fsm_42_1 = 1;
  localparam _mystream_b10_source_fsm_42_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_b10_source_fsm_42 <= _mystream_b10_source_fsm_42_init;
    end else begin
      case(_mystream_b10_source_fsm_42)
        _mystream_b10_source_fsm_42_init: begin
          if(_mystream_source_start && _mystream_b10_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_b10_source_fsm_42 <= _mystream_b10_source_fsm_42_1;
          end 
        end
        _mystream_b10_source_fsm_42_1: begin
          if(_mystream_stream_oready) begin
            _mystream_b10_source_fsm_42 <= _mystream_b10_source_fsm_42_2;
          end 
        end
        _mystream_b10_source_fsm_42_2: begin
          if((_mystream_b10_source_count == 1) && _mystream_stream_oready) begin
            _mystream_b10_source_fsm_42 <= _mystream_b10_source_fsm_42_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_b10_source_fsm_42 <= _mystream_b10_source_fsm_42_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_b11_source_fsm_43_1 = 1;
  localparam _mystream_b11_source_fsm_43_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_b11_source_fsm_43 <= _mystream_b11_source_fsm_43_init;
    end else begin
      case(_mystream_b11_source_fsm_43)
        _mystream_b11_source_fsm_43_init: begin
          if(_mystream_source_start && _mystream_b11_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_b11_source_fsm_43 <= _mystream_b11_source_fsm_43_1;
          end 
        end
        _mystream_b11_source_fsm_43_1: begin
          if(_mystream_stream_oready) begin
            _mystream_b11_source_fsm_43 <= _mystream_b11_source_fsm_43_2;
          end 
        end
        _mystream_b11_source_fsm_43_2: begin
          if((_mystream_b11_source_count == 1) && _mystream_stream_oready) begin
            _mystream_b11_source_fsm_43 <= _mystream_b11_source_fsm_43_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_b11_source_fsm_43 <= _mystream_b11_source_fsm_43_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_b12_source_fsm_44_1 = 1;
  localparam _mystream_b12_source_fsm_44_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_b12_source_fsm_44 <= _mystream_b12_source_fsm_44_init;
    end else begin
      case(_mystream_b12_source_fsm_44)
        _mystream_b12_source_fsm_44_init: begin
          if(_mystream_source_start && _mystream_b12_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_b12_source_fsm_44 <= _mystream_b12_source_fsm_44_1;
          end 
        end
        _mystream_b12_source_fsm_44_1: begin
          if(_mystream_stream_oready) begin
            _mystream_b12_source_fsm_44 <= _mystream_b12_source_fsm_44_2;
          end 
        end
        _mystream_b12_source_fsm_44_2: begin
          if((_mystream_b12_source_count == 1) && _mystream_stream_oready) begin
            _mystream_b12_source_fsm_44 <= _mystream_b12_source_fsm_44_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_b12_source_fsm_44 <= _mystream_b12_source_fsm_44_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_b13_source_fsm_45_1 = 1;
  localparam _mystream_b13_source_fsm_45_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_b13_source_fsm_45 <= _mystream_b13_source_fsm_45_init;
    end else begin
      case(_mystream_b13_source_fsm_45)
        _mystream_b13_source_fsm_45_init: begin
          if(_mystream_source_start && _mystream_b13_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_b13_source_fsm_45 <= _mystream_b13_source_fsm_45_1;
          end 
        end
        _mystream_b13_source_fsm_45_1: begin
          if(_mystream_stream_oready) begin
            _mystream_b13_source_fsm_45 <= _mystream_b13_source_fsm_45_2;
          end 
        end
        _mystream_b13_source_fsm_45_2: begin
          if((_mystream_b13_source_count == 1) && _mystream_stream_oready) begin
            _mystream_b13_source_fsm_45 <= _mystream_b13_source_fsm_45_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_b13_source_fsm_45 <= _mystream_b13_source_fsm_45_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_b14_source_fsm_46_1 = 1;
  localparam _mystream_b14_source_fsm_46_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_b14_source_fsm_46 <= _mystream_b14_source_fsm_46_init;
    end else begin
      case(_mystream_b14_source_fsm_46)
        _mystream_b14_source_fsm_46_init: begin
          if(_mystream_source_start && _mystream_b14_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_b14_source_fsm_46 <= _mystream_b14_source_fsm_46_1;
          end 
        end
        _mystream_b14_source_fsm_46_1: begin
          if(_mystream_stream_oready) begin
            _mystream_b14_source_fsm_46 <= _mystream_b14_source_fsm_46_2;
          end 
        end
        _mystream_b14_source_fsm_46_2: begin
          if((_mystream_b14_source_count == 1) && _mystream_stream_oready) begin
            _mystream_b14_source_fsm_46 <= _mystream_b14_source_fsm_46_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_b14_source_fsm_46 <= _mystream_b14_source_fsm_46_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_b15_source_fsm_47_1 = 1;
  localparam _mystream_b15_source_fsm_47_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_b15_source_fsm_47 <= _mystream_b15_source_fsm_47_init;
    end else begin
      case(_mystream_b15_source_fsm_47)
        _mystream_b15_source_fsm_47_init: begin
          if(_mystream_source_start && _mystream_b15_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_b15_source_fsm_47 <= _mystream_b15_source_fsm_47_1;
          end 
        end
        _mystream_b15_source_fsm_47_1: begin
          if(_mystream_stream_oready) begin
            _mystream_b15_source_fsm_47 <= _mystream_b15_source_fsm_47_2;
          end 
        end
        _mystream_b15_source_fsm_47_2: begin
          if((_mystream_b15_source_count == 1) && _mystream_stream_oready) begin
            _mystream_b15_source_fsm_47 <= _mystream_b15_source_fsm_47_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_b15_source_fsm_47 <= _mystream_b15_source_fsm_47_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_b16_source_fsm_48_1 = 1;
  localparam _mystream_b16_source_fsm_48_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_b16_source_fsm_48 <= _mystream_b16_source_fsm_48_init;
    end else begin
      case(_mystream_b16_source_fsm_48)
        _mystream_b16_source_fsm_48_init: begin
          if(_mystream_source_start && _mystream_b16_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_b16_source_fsm_48 <= _mystream_b16_source_fsm_48_1;
          end 
        end
        _mystream_b16_source_fsm_48_1: begin
          if(_mystream_stream_oready) begin
            _mystream_b16_source_fsm_48 <= _mystream_b16_source_fsm_48_2;
          end 
        end
        _mystream_b16_source_fsm_48_2: begin
          if((_mystream_b16_source_count == 1) && _mystream_stream_oready) begin
            _mystream_b16_source_fsm_48 <= _mystream_b16_source_fsm_48_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_b16_source_fsm_48 <= _mystream_b16_source_fsm_48_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_b17_source_fsm_49_1 = 1;
  localparam _mystream_b17_source_fsm_49_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_b17_source_fsm_49 <= _mystream_b17_source_fsm_49_init;
    end else begin
      case(_mystream_b17_source_fsm_49)
        _mystream_b17_source_fsm_49_init: begin
          if(_mystream_source_start && _mystream_b17_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_b17_source_fsm_49 <= _mystream_b17_source_fsm_49_1;
          end 
        end
        _mystream_b17_source_fsm_49_1: begin
          if(_mystream_stream_oready) begin
            _mystream_b17_source_fsm_49 <= _mystream_b17_source_fsm_49_2;
          end 
        end
        _mystream_b17_source_fsm_49_2: begin
          if((_mystream_b17_source_count == 1) && _mystream_stream_oready) begin
            _mystream_b17_source_fsm_49 <= _mystream_b17_source_fsm_49_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_b17_source_fsm_49 <= _mystream_b17_source_fsm_49_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_b18_source_fsm_50_1 = 1;
  localparam _mystream_b18_source_fsm_50_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_b18_source_fsm_50 <= _mystream_b18_source_fsm_50_init;
    end else begin
      case(_mystream_b18_source_fsm_50)
        _mystream_b18_source_fsm_50_init: begin
          if(_mystream_source_start && _mystream_b18_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_b18_source_fsm_50 <= _mystream_b18_source_fsm_50_1;
          end 
        end
        _mystream_b18_source_fsm_50_1: begin
          if(_mystream_stream_oready) begin
            _mystream_b18_source_fsm_50 <= _mystream_b18_source_fsm_50_2;
          end 
        end
        _mystream_b18_source_fsm_50_2: begin
          if((_mystream_b18_source_count == 1) && _mystream_stream_oready) begin
            _mystream_b18_source_fsm_50 <= _mystream_b18_source_fsm_50_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_b18_source_fsm_50 <= _mystream_b18_source_fsm_50_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_b19_source_fsm_51_1 = 1;
  localparam _mystream_b19_source_fsm_51_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_b19_source_fsm_51 <= _mystream_b19_source_fsm_51_init;
    end else begin
      case(_mystream_b19_source_fsm_51)
        _mystream_b19_source_fsm_51_init: begin
          if(_mystream_source_start && _mystream_b19_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_b19_source_fsm_51 <= _mystream_b19_source_fsm_51_1;
          end 
        end
        _mystream_b19_source_fsm_51_1: begin
          if(_mystream_stream_oready) begin
            _mystream_b19_source_fsm_51 <= _mystream_b19_source_fsm_51_2;
          end 
        end
        _mystream_b19_source_fsm_51_2: begin
          if((_mystream_b19_source_count == 1) && _mystream_stream_oready) begin
            _mystream_b19_source_fsm_51 <= _mystream_b19_source_fsm_51_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_b19_source_fsm_51 <= _mystream_b19_source_fsm_51_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_b20_source_fsm_52_1 = 1;
  localparam _mystream_b20_source_fsm_52_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_b20_source_fsm_52 <= _mystream_b20_source_fsm_52_init;
    end else begin
      case(_mystream_b20_source_fsm_52)
        _mystream_b20_source_fsm_52_init: begin
          if(_mystream_source_start && _mystream_b20_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_b20_source_fsm_52 <= _mystream_b20_source_fsm_52_1;
          end 
        end
        _mystream_b20_source_fsm_52_1: begin
          if(_mystream_stream_oready) begin
            _mystream_b20_source_fsm_52 <= _mystream_b20_source_fsm_52_2;
          end 
        end
        _mystream_b20_source_fsm_52_2: begin
          if((_mystream_b20_source_count == 1) && _mystream_stream_oready) begin
            _mystream_b20_source_fsm_52 <= _mystream_b20_source_fsm_52_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_b20_source_fsm_52 <= _mystream_b20_source_fsm_52_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_b21_source_fsm_53_1 = 1;
  localparam _mystream_b21_source_fsm_53_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_b21_source_fsm_53 <= _mystream_b21_source_fsm_53_init;
    end else begin
      case(_mystream_b21_source_fsm_53)
        _mystream_b21_source_fsm_53_init: begin
          if(_mystream_source_start && _mystream_b21_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_b21_source_fsm_53 <= _mystream_b21_source_fsm_53_1;
          end 
        end
        _mystream_b21_source_fsm_53_1: begin
          if(_mystream_stream_oready) begin
            _mystream_b21_source_fsm_53 <= _mystream_b21_source_fsm_53_2;
          end 
        end
        _mystream_b21_source_fsm_53_2: begin
          if((_mystream_b21_source_count == 1) && _mystream_stream_oready) begin
            _mystream_b21_source_fsm_53 <= _mystream_b21_source_fsm_53_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_b21_source_fsm_53 <= _mystream_b21_source_fsm_53_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_b22_source_fsm_54_1 = 1;
  localparam _mystream_b22_source_fsm_54_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_b22_source_fsm_54 <= _mystream_b22_source_fsm_54_init;
    end else begin
      case(_mystream_b22_source_fsm_54)
        _mystream_b22_source_fsm_54_init: begin
          if(_mystream_source_start && _mystream_b22_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_b22_source_fsm_54 <= _mystream_b22_source_fsm_54_1;
          end 
        end
        _mystream_b22_source_fsm_54_1: begin
          if(_mystream_stream_oready) begin
            _mystream_b22_source_fsm_54 <= _mystream_b22_source_fsm_54_2;
          end 
        end
        _mystream_b22_source_fsm_54_2: begin
          if((_mystream_b22_source_count == 1) && _mystream_stream_oready) begin
            _mystream_b22_source_fsm_54 <= _mystream_b22_source_fsm_54_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_b22_source_fsm_54 <= _mystream_b22_source_fsm_54_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_b23_source_fsm_55_1 = 1;
  localparam _mystream_b23_source_fsm_55_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_b23_source_fsm_55 <= _mystream_b23_source_fsm_55_init;
    end else begin
      case(_mystream_b23_source_fsm_55)
        _mystream_b23_source_fsm_55_init: begin
          if(_mystream_source_start && _mystream_b23_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_b23_source_fsm_55 <= _mystream_b23_source_fsm_55_1;
          end 
        end
        _mystream_b23_source_fsm_55_1: begin
          if(_mystream_stream_oready) begin
            _mystream_b23_source_fsm_55 <= _mystream_b23_source_fsm_55_2;
          end 
        end
        _mystream_b23_source_fsm_55_2: begin
          if((_mystream_b23_source_count == 1) && _mystream_stream_oready) begin
            _mystream_b23_source_fsm_55 <= _mystream_b23_source_fsm_55_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_b23_source_fsm_55 <= _mystream_b23_source_fsm_55_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_b24_source_fsm_56_1 = 1;
  localparam _mystream_b24_source_fsm_56_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_b24_source_fsm_56 <= _mystream_b24_source_fsm_56_init;
    end else begin
      case(_mystream_b24_source_fsm_56)
        _mystream_b24_source_fsm_56_init: begin
          if(_mystream_source_start && _mystream_b24_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_b24_source_fsm_56 <= _mystream_b24_source_fsm_56_1;
          end 
        end
        _mystream_b24_source_fsm_56_1: begin
          if(_mystream_stream_oready) begin
            _mystream_b24_source_fsm_56 <= _mystream_b24_source_fsm_56_2;
          end 
        end
        _mystream_b24_source_fsm_56_2: begin
          if((_mystream_b24_source_count == 1) && _mystream_stream_oready) begin
            _mystream_b24_source_fsm_56 <= _mystream_b24_source_fsm_56_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_b24_source_fsm_56 <= _mystream_b24_source_fsm_56_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_b25_source_fsm_57_1 = 1;
  localparam _mystream_b25_source_fsm_57_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_b25_source_fsm_57 <= _mystream_b25_source_fsm_57_init;
    end else begin
      case(_mystream_b25_source_fsm_57)
        _mystream_b25_source_fsm_57_init: begin
          if(_mystream_source_start && _mystream_b25_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_b25_source_fsm_57 <= _mystream_b25_source_fsm_57_1;
          end 
        end
        _mystream_b25_source_fsm_57_1: begin
          if(_mystream_stream_oready) begin
            _mystream_b25_source_fsm_57 <= _mystream_b25_source_fsm_57_2;
          end 
        end
        _mystream_b25_source_fsm_57_2: begin
          if((_mystream_b25_source_count == 1) && _mystream_stream_oready) begin
            _mystream_b25_source_fsm_57 <= _mystream_b25_source_fsm_57_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_b25_source_fsm_57 <= _mystream_b25_source_fsm_57_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_b26_source_fsm_58_1 = 1;
  localparam _mystream_b26_source_fsm_58_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_b26_source_fsm_58 <= _mystream_b26_source_fsm_58_init;
    end else begin
      case(_mystream_b26_source_fsm_58)
        _mystream_b26_source_fsm_58_init: begin
          if(_mystream_source_start && _mystream_b26_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_b26_source_fsm_58 <= _mystream_b26_source_fsm_58_1;
          end 
        end
        _mystream_b26_source_fsm_58_1: begin
          if(_mystream_stream_oready) begin
            _mystream_b26_source_fsm_58 <= _mystream_b26_source_fsm_58_2;
          end 
        end
        _mystream_b26_source_fsm_58_2: begin
          if((_mystream_b26_source_count == 1) && _mystream_stream_oready) begin
            _mystream_b26_source_fsm_58 <= _mystream_b26_source_fsm_58_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_b26_source_fsm_58 <= _mystream_b26_source_fsm_58_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_b27_source_fsm_59_1 = 1;
  localparam _mystream_b27_source_fsm_59_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_b27_source_fsm_59 <= _mystream_b27_source_fsm_59_init;
    end else begin
      case(_mystream_b27_source_fsm_59)
        _mystream_b27_source_fsm_59_init: begin
          if(_mystream_source_start && _mystream_b27_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_b27_source_fsm_59 <= _mystream_b27_source_fsm_59_1;
          end 
        end
        _mystream_b27_source_fsm_59_1: begin
          if(_mystream_stream_oready) begin
            _mystream_b27_source_fsm_59 <= _mystream_b27_source_fsm_59_2;
          end 
        end
        _mystream_b27_source_fsm_59_2: begin
          if((_mystream_b27_source_count == 1) && _mystream_stream_oready) begin
            _mystream_b27_source_fsm_59 <= _mystream_b27_source_fsm_59_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_b27_source_fsm_59 <= _mystream_b27_source_fsm_59_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_b28_source_fsm_60_1 = 1;
  localparam _mystream_b28_source_fsm_60_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_b28_source_fsm_60 <= _mystream_b28_source_fsm_60_init;
    end else begin
      case(_mystream_b28_source_fsm_60)
        _mystream_b28_source_fsm_60_init: begin
          if(_mystream_source_start && _mystream_b28_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_b28_source_fsm_60 <= _mystream_b28_source_fsm_60_1;
          end 
        end
        _mystream_b28_source_fsm_60_1: begin
          if(_mystream_stream_oready) begin
            _mystream_b28_source_fsm_60 <= _mystream_b28_source_fsm_60_2;
          end 
        end
        _mystream_b28_source_fsm_60_2: begin
          if((_mystream_b28_source_count == 1) && _mystream_stream_oready) begin
            _mystream_b28_source_fsm_60 <= _mystream_b28_source_fsm_60_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_b28_source_fsm_60 <= _mystream_b28_source_fsm_60_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_b29_source_fsm_61_1 = 1;
  localparam _mystream_b29_source_fsm_61_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_b29_source_fsm_61 <= _mystream_b29_source_fsm_61_init;
    end else begin
      case(_mystream_b29_source_fsm_61)
        _mystream_b29_source_fsm_61_init: begin
          if(_mystream_source_start && _mystream_b29_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_b29_source_fsm_61 <= _mystream_b29_source_fsm_61_1;
          end 
        end
        _mystream_b29_source_fsm_61_1: begin
          if(_mystream_stream_oready) begin
            _mystream_b29_source_fsm_61 <= _mystream_b29_source_fsm_61_2;
          end 
        end
        _mystream_b29_source_fsm_61_2: begin
          if((_mystream_b29_source_count == 1) && _mystream_stream_oready) begin
            _mystream_b29_source_fsm_61 <= _mystream_b29_source_fsm_61_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_b29_source_fsm_61 <= _mystream_b29_source_fsm_61_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_b30_source_fsm_62_1 = 1;
  localparam _mystream_b30_source_fsm_62_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_b30_source_fsm_62 <= _mystream_b30_source_fsm_62_init;
    end else begin
      case(_mystream_b30_source_fsm_62)
        _mystream_b30_source_fsm_62_init: begin
          if(_mystream_source_start && _mystream_b30_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_b30_source_fsm_62 <= _mystream_b30_source_fsm_62_1;
          end 
        end
        _mystream_b30_source_fsm_62_1: begin
          if(_mystream_stream_oready) begin
            _mystream_b30_source_fsm_62 <= _mystream_b30_source_fsm_62_2;
          end 
        end
        _mystream_b30_source_fsm_62_2: begin
          if((_mystream_b30_source_count == 1) && _mystream_stream_oready) begin
            _mystream_b30_source_fsm_62 <= _mystream_b30_source_fsm_62_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_b30_source_fsm_62 <= _mystream_b30_source_fsm_62_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_b31_source_fsm_63_1 = 1;
  localparam _mystream_b31_source_fsm_63_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_b31_source_fsm_63 <= _mystream_b31_source_fsm_63_init;
    end else begin
      case(_mystream_b31_source_fsm_63)
        _mystream_b31_source_fsm_63_init: begin
          if(_mystream_source_start && _mystream_b31_source_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_b31_source_fsm_63 <= _mystream_b31_source_fsm_63_1;
          end 
        end
        _mystream_b31_source_fsm_63_1: begin
          if(_mystream_stream_oready) begin
            _mystream_b31_source_fsm_63 <= _mystream_b31_source_fsm_63_2;
          end 
        end
        _mystream_b31_source_fsm_63_2: begin
          if((_mystream_b31_source_count == 1) && _mystream_stream_oready) begin
            _mystream_b31_source_fsm_63 <= _mystream_b31_source_fsm_63_init;
          end 
          if(_mystream_source_stop && _mystream_stream_oready) begin
            _mystream_b31_source_fsm_63 <= _mystream_b31_source_fsm_63_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_sum_vec0_sink_fsm_64_1 = 1;
  localparam _mystream_sum_vec0_sink_fsm_64_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_sum_vec0_sink_fsm_64 <= _mystream_sum_vec0_sink_fsm_64_init;
    end else begin
      case(_mystream_sum_vec0_sink_fsm_64)
        _mystream_sum_vec0_sink_fsm_64_init: begin
          if(_mystream_sink_start && _mystream_sum_vec0_sink_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_sum_vec0_sink_fsm_64 <= _mystream_sum_vec0_sink_fsm_64_1;
          end 
        end
        _mystream_sum_vec0_sink_fsm_64_1: begin
          if(_mystream_stream_oready) begin
            _mystream_sum_vec0_sink_fsm_64 <= _mystream_sum_vec0_sink_fsm_64_2;
          end 
        end
        _mystream_sum_vec0_sink_fsm_64_2: begin
          if((_mystream_sum_vec0_sink_count == 1) && _mystream_stream_oready) begin
            _mystream_sum_vec0_sink_fsm_64 <= _mystream_sum_vec0_sink_fsm_64_init;
          end 
          if(_mystream_sink_stop && _mystream_stream_oready) begin
            _mystream_sum_vec0_sink_fsm_64 <= _mystream_sum_vec0_sink_fsm_64_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_sum_vec1_sink_fsm_65_1 = 1;
  localparam _mystream_sum_vec1_sink_fsm_65_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_sum_vec1_sink_fsm_65 <= _mystream_sum_vec1_sink_fsm_65_init;
    end else begin
      case(_mystream_sum_vec1_sink_fsm_65)
        _mystream_sum_vec1_sink_fsm_65_init: begin
          if(_mystream_sink_start && _mystream_sum_vec1_sink_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_sum_vec1_sink_fsm_65 <= _mystream_sum_vec1_sink_fsm_65_1;
          end 
        end
        _mystream_sum_vec1_sink_fsm_65_1: begin
          if(_mystream_stream_oready) begin
            _mystream_sum_vec1_sink_fsm_65 <= _mystream_sum_vec1_sink_fsm_65_2;
          end 
        end
        _mystream_sum_vec1_sink_fsm_65_2: begin
          if((_mystream_sum_vec1_sink_count == 1) && _mystream_stream_oready) begin
            _mystream_sum_vec1_sink_fsm_65 <= _mystream_sum_vec1_sink_fsm_65_init;
          end 
          if(_mystream_sink_stop && _mystream_stream_oready) begin
            _mystream_sum_vec1_sink_fsm_65 <= _mystream_sum_vec1_sink_fsm_65_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_sum_vec2_sink_fsm_66_1 = 1;
  localparam _mystream_sum_vec2_sink_fsm_66_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_sum_vec2_sink_fsm_66 <= _mystream_sum_vec2_sink_fsm_66_init;
    end else begin
      case(_mystream_sum_vec2_sink_fsm_66)
        _mystream_sum_vec2_sink_fsm_66_init: begin
          if(_mystream_sink_start && _mystream_sum_vec2_sink_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_sum_vec2_sink_fsm_66 <= _mystream_sum_vec2_sink_fsm_66_1;
          end 
        end
        _mystream_sum_vec2_sink_fsm_66_1: begin
          if(_mystream_stream_oready) begin
            _mystream_sum_vec2_sink_fsm_66 <= _mystream_sum_vec2_sink_fsm_66_2;
          end 
        end
        _mystream_sum_vec2_sink_fsm_66_2: begin
          if((_mystream_sum_vec2_sink_count == 1) && _mystream_stream_oready) begin
            _mystream_sum_vec2_sink_fsm_66 <= _mystream_sum_vec2_sink_fsm_66_init;
          end 
          if(_mystream_sink_stop && _mystream_stream_oready) begin
            _mystream_sum_vec2_sink_fsm_66 <= _mystream_sum_vec2_sink_fsm_66_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_sum_vec3_sink_fsm_67_1 = 1;
  localparam _mystream_sum_vec3_sink_fsm_67_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_sum_vec3_sink_fsm_67 <= _mystream_sum_vec3_sink_fsm_67_init;
    end else begin
      case(_mystream_sum_vec3_sink_fsm_67)
        _mystream_sum_vec3_sink_fsm_67_init: begin
          if(_mystream_sink_start && _mystream_sum_vec3_sink_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_sum_vec3_sink_fsm_67 <= _mystream_sum_vec3_sink_fsm_67_1;
          end 
        end
        _mystream_sum_vec3_sink_fsm_67_1: begin
          if(_mystream_stream_oready) begin
            _mystream_sum_vec3_sink_fsm_67 <= _mystream_sum_vec3_sink_fsm_67_2;
          end 
        end
        _mystream_sum_vec3_sink_fsm_67_2: begin
          if((_mystream_sum_vec3_sink_count == 1) && _mystream_stream_oready) begin
            _mystream_sum_vec3_sink_fsm_67 <= _mystream_sum_vec3_sink_fsm_67_init;
          end 
          if(_mystream_sink_stop && _mystream_stream_oready) begin
            _mystream_sum_vec3_sink_fsm_67 <= _mystream_sum_vec3_sink_fsm_67_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_sum_vec4_sink_fsm_68_1 = 1;
  localparam _mystream_sum_vec4_sink_fsm_68_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_sum_vec4_sink_fsm_68 <= _mystream_sum_vec4_sink_fsm_68_init;
    end else begin
      case(_mystream_sum_vec4_sink_fsm_68)
        _mystream_sum_vec4_sink_fsm_68_init: begin
          if(_mystream_sink_start && _mystream_sum_vec4_sink_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_sum_vec4_sink_fsm_68 <= _mystream_sum_vec4_sink_fsm_68_1;
          end 
        end
        _mystream_sum_vec4_sink_fsm_68_1: begin
          if(_mystream_stream_oready) begin
            _mystream_sum_vec4_sink_fsm_68 <= _mystream_sum_vec4_sink_fsm_68_2;
          end 
        end
        _mystream_sum_vec4_sink_fsm_68_2: begin
          if((_mystream_sum_vec4_sink_count == 1) && _mystream_stream_oready) begin
            _mystream_sum_vec4_sink_fsm_68 <= _mystream_sum_vec4_sink_fsm_68_init;
          end 
          if(_mystream_sink_stop && _mystream_stream_oready) begin
            _mystream_sum_vec4_sink_fsm_68 <= _mystream_sum_vec4_sink_fsm_68_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_sum_vec5_sink_fsm_69_1 = 1;
  localparam _mystream_sum_vec5_sink_fsm_69_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_sum_vec5_sink_fsm_69 <= _mystream_sum_vec5_sink_fsm_69_init;
    end else begin
      case(_mystream_sum_vec5_sink_fsm_69)
        _mystream_sum_vec5_sink_fsm_69_init: begin
          if(_mystream_sink_start && _mystream_sum_vec5_sink_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_sum_vec5_sink_fsm_69 <= _mystream_sum_vec5_sink_fsm_69_1;
          end 
        end
        _mystream_sum_vec5_sink_fsm_69_1: begin
          if(_mystream_stream_oready) begin
            _mystream_sum_vec5_sink_fsm_69 <= _mystream_sum_vec5_sink_fsm_69_2;
          end 
        end
        _mystream_sum_vec5_sink_fsm_69_2: begin
          if((_mystream_sum_vec5_sink_count == 1) && _mystream_stream_oready) begin
            _mystream_sum_vec5_sink_fsm_69 <= _mystream_sum_vec5_sink_fsm_69_init;
          end 
          if(_mystream_sink_stop && _mystream_stream_oready) begin
            _mystream_sum_vec5_sink_fsm_69 <= _mystream_sum_vec5_sink_fsm_69_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_sum_vec6_sink_fsm_70_1 = 1;
  localparam _mystream_sum_vec6_sink_fsm_70_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_sum_vec6_sink_fsm_70 <= _mystream_sum_vec6_sink_fsm_70_init;
    end else begin
      case(_mystream_sum_vec6_sink_fsm_70)
        _mystream_sum_vec6_sink_fsm_70_init: begin
          if(_mystream_sink_start && _mystream_sum_vec6_sink_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_sum_vec6_sink_fsm_70 <= _mystream_sum_vec6_sink_fsm_70_1;
          end 
        end
        _mystream_sum_vec6_sink_fsm_70_1: begin
          if(_mystream_stream_oready) begin
            _mystream_sum_vec6_sink_fsm_70 <= _mystream_sum_vec6_sink_fsm_70_2;
          end 
        end
        _mystream_sum_vec6_sink_fsm_70_2: begin
          if((_mystream_sum_vec6_sink_count == 1) && _mystream_stream_oready) begin
            _mystream_sum_vec6_sink_fsm_70 <= _mystream_sum_vec6_sink_fsm_70_init;
          end 
          if(_mystream_sink_stop && _mystream_stream_oready) begin
            _mystream_sum_vec6_sink_fsm_70 <= _mystream_sum_vec6_sink_fsm_70_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_sum_vec7_sink_fsm_71_1 = 1;
  localparam _mystream_sum_vec7_sink_fsm_71_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_sum_vec7_sink_fsm_71 <= _mystream_sum_vec7_sink_fsm_71_init;
    end else begin
      case(_mystream_sum_vec7_sink_fsm_71)
        _mystream_sum_vec7_sink_fsm_71_init: begin
          if(_mystream_sink_start && _mystream_sum_vec7_sink_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_sum_vec7_sink_fsm_71 <= _mystream_sum_vec7_sink_fsm_71_1;
          end 
        end
        _mystream_sum_vec7_sink_fsm_71_1: begin
          if(_mystream_stream_oready) begin
            _mystream_sum_vec7_sink_fsm_71 <= _mystream_sum_vec7_sink_fsm_71_2;
          end 
        end
        _mystream_sum_vec7_sink_fsm_71_2: begin
          if((_mystream_sum_vec7_sink_count == 1) && _mystream_stream_oready) begin
            _mystream_sum_vec7_sink_fsm_71 <= _mystream_sum_vec7_sink_fsm_71_init;
          end 
          if(_mystream_sink_stop && _mystream_stream_oready) begin
            _mystream_sum_vec7_sink_fsm_71 <= _mystream_sum_vec7_sink_fsm_71_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_sum_vec8_sink_fsm_72_1 = 1;
  localparam _mystream_sum_vec8_sink_fsm_72_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_sum_vec8_sink_fsm_72 <= _mystream_sum_vec8_sink_fsm_72_init;
    end else begin
      case(_mystream_sum_vec8_sink_fsm_72)
        _mystream_sum_vec8_sink_fsm_72_init: begin
          if(_mystream_sink_start && _mystream_sum_vec8_sink_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_sum_vec8_sink_fsm_72 <= _mystream_sum_vec8_sink_fsm_72_1;
          end 
        end
        _mystream_sum_vec8_sink_fsm_72_1: begin
          if(_mystream_stream_oready) begin
            _mystream_sum_vec8_sink_fsm_72 <= _mystream_sum_vec8_sink_fsm_72_2;
          end 
        end
        _mystream_sum_vec8_sink_fsm_72_2: begin
          if((_mystream_sum_vec8_sink_count == 1) && _mystream_stream_oready) begin
            _mystream_sum_vec8_sink_fsm_72 <= _mystream_sum_vec8_sink_fsm_72_init;
          end 
          if(_mystream_sink_stop && _mystream_stream_oready) begin
            _mystream_sum_vec8_sink_fsm_72 <= _mystream_sum_vec8_sink_fsm_72_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_sum_vec9_sink_fsm_73_1 = 1;
  localparam _mystream_sum_vec9_sink_fsm_73_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_sum_vec9_sink_fsm_73 <= _mystream_sum_vec9_sink_fsm_73_init;
    end else begin
      case(_mystream_sum_vec9_sink_fsm_73)
        _mystream_sum_vec9_sink_fsm_73_init: begin
          if(_mystream_sink_start && _mystream_sum_vec9_sink_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_sum_vec9_sink_fsm_73 <= _mystream_sum_vec9_sink_fsm_73_1;
          end 
        end
        _mystream_sum_vec9_sink_fsm_73_1: begin
          if(_mystream_stream_oready) begin
            _mystream_sum_vec9_sink_fsm_73 <= _mystream_sum_vec9_sink_fsm_73_2;
          end 
        end
        _mystream_sum_vec9_sink_fsm_73_2: begin
          if((_mystream_sum_vec9_sink_count == 1) && _mystream_stream_oready) begin
            _mystream_sum_vec9_sink_fsm_73 <= _mystream_sum_vec9_sink_fsm_73_init;
          end 
          if(_mystream_sink_stop && _mystream_stream_oready) begin
            _mystream_sum_vec9_sink_fsm_73 <= _mystream_sum_vec9_sink_fsm_73_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_sum_vec10_sink_fsm_74_1 = 1;
  localparam _mystream_sum_vec10_sink_fsm_74_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_sum_vec10_sink_fsm_74 <= _mystream_sum_vec10_sink_fsm_74_init;
    end else begin
      case(_mystream_sum_vec10_sink_fsm_74)
        _mystream_sum_vec10_sink_fsm_74_init: begin
          if(_mystream_sink_start && _mystream_sum_vec10_sink_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_sum_vec10_sink_fsm_74 <= _mystream_sum_vec10_sink_fsm_74_1;
          end 
        end
        _mystream_sum_vec10_sink_fsm_74_1: begin
          if(_mystream_stream_oready) begin
            _mystream_sum_vec10_sink_fsm_74 <= _mystream_sum_vec10_sink_fsm_74_2;
          end 
        end
        _mystream_sum_vec10_sink_fsm_74_2: begin
          if((_mystream_sum_vec10_sink_count == 1) && _mystream_stream_oready) begin
            _mystream_sum_vec10_sink_fsm_74 <= _mystream_sum_vec10_sink_fsm_74_init;
          end 
          if(_mystream_sink_stop && _mystream_stream_oready) begin
            _mystream_sum_vec10_sink_fsm_74 <= _mystream_sum_vec10_sink_fsm_74_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_sum_vec11_sink_fsm_75_1 = 1;
  localparam _mystream_sum_vec11_sink_fsm_75_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_sum_vec11_sink_fsm_75 <= _mystream_sum_vec11_sink_fsm_75_init;
    end else begin
      case(_mystream_sum_vec11_sink_fsm_75)
        _mystream_sum_vec11_sink_fsm_75_init: begin
          if(_mystream_sink_start && _mystream_sum_vec11_sink_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_sum_vec11_sink_fsm_75 <= _mystream_sum_vec11_sink_fsm_75_1;
          end 
        end
        _mystream_sum_vec11_sink_fsm_75_1: begin
          if(_mystream_stream_oready) begin
            _mystream_sum_vec11_sink_fsm_75 <= _mystream_sum_vec11_sink_fsm_75_2;
          end 
        end
        _mystream_sum_vec11_sink_fsm_75_2: begin
          if((_mystream_sum_vec11_sink_count == 1) && _mystream_stream_oready) begin
            _mystream_sum_vec11_sink_fsm_75 <= _mystream_sum_vec11_sink_fsm_75_init;
          end 
          if(_mystream_sink_stop && _mystream_stream_oready) begin
            _mystream_sum_vec11_sink_fsm_75 <= _mystream_sum_vec11_sink_fsm_75_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_sum_vec12_sink_fsm_76_1 = 1;
  localparam _mystream_sum_vec12_sink_fsm_76_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_sum_vec12_sink_fsm_76 <= _mystream_sum_vec12_sink_fsm_76_init;
    end else begin
      case(_mystream_sum_vec12_sink_fsm_76)
        _mystream_sum_vec12_sink_fsm_76_init: begin
          if(_mystream_sink_start && _mystream_sum_vec12_sink_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_sum_vec12_sink_fsm_76 <= _mystream_sum_vec12_sink_fsm_76_1;
          end 
        end
        _mystream_sum_vec12_sink_fsm_76_1: begin
          if(_mystream_stream_oready) begin
            _mystream_sum_vec12_sink_fsm_76 <= _mystream_sum_vec12_sink_fsm_76_2;
          end 
        end
        _mystream_sum_vec12_sink_fsm_76_2: begin
          if((_mystream_sum_vec12_sink_count == 1) && _mystream_stream_oready) begin
            _mystream_sum_vec12_sink_fsm_76 <= _mystream_sum_vec12_sink_fsm_76_init;
          end 
          if(_mystream_sink_stop && _mystream_stream_oready) begin
            _mystream_sum_vec12_sink_fsm_76 <= _mystream_sum_vec12_sink_fsm_76_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_sum_vec13_sink_fsm_77_1 = 1;
  localparam _mystream_sum_vec13_sink_fsm_77_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_sum_vec13_sink_fsm_77 <= _mystream_sum_vec13_sink_fsm_77_init;
    end else begin
      case(_mystream_sum_vec13_sink_fsm_77)
        _mystream_sum_vec13_sink_fsm_77_init: begin
          if(_mystream_sink_start && _mystream_sum_vec13_sink_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_sum_vec13_sink_fsm_77 <= _mystream_sum_vec13_sink_fsm_77_1;
          end 
        end
        _mystream_sum_vec13_sink_fsm_77_1: begin
          if(_mystream_stream_oready) begin
            _mystream_sum_vec13_sink_fsm_77 <= _mystream_sum_vec13_sink_fsm_77_2;
          end 
        end
        _mystream_sum_vec13_sink_fsm_77_2: begin
          if((_mystream_sum_vec13_sink_count == 1) && _mystream_stream_oready) begin
            _mystream_sum_vec13_sink_fsm_77 <= _mystream_sum_vec13_sink_fsm_77_init;
          end 
          if(_mystream_sink_stop && _mystream_stream_oready) begin
            _mystream_sum_vec13_sink_fsm_77 <= _mystream_sum_vec13_sink_fsm_77_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_sum_vec14_sink_fsm_78_1 = 1;
  localparam _mystream_sum_vec14_sink_fsm_78_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_sum_vec14_sink_fsm_78 <= _mystream_sum_vec14_sink_fsm_78_init;
    end else begin
      case(_mystream_sum_vec14_sink_fsm_78)
        _mystream_sum_vec14_sink_fsm_78_init: begin
          if(_mystream_sink_start && _mystream_sum_vec14_sink_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_sum_vec14_sink_fsm_78 <= _mystream_sum_vec14_sink_fsm_78_1;
          end 
        end
        _mystream_sum_vec14_sink_fsm_78_1: begin
          if(_mystream_stream_oready) begin
            _mystream_sum_vec14_sink_fsm_78 <= _mystream_sum_vec14_sink_fsm_78_2;
          end 
        end
        _mystream_sum_vec14_sink_fsm_78_2: begin
          if((_mystream_sum_vec14_sink_count == 1) && _mystream_stream_oready) begin
            _mystream_sum_vec14_sink_fsm_78 <= _mystream_sum_vec14_sink_fsm_78_init;
          end 
          if(_mystream_sink_stop && _mystream_stream_oready) begin
            _mystream_sum_vec14_sink_fsm_78 <= _mystream_sum_vec14_sink_fsm_78_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_sum_vec15_sink_fsm_79_1 = 1;
  localparam _mystream_sum_vec15_sink_fsm_79_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_sum_vec15_sink_fsm_79 <= _mystream_sum_vec15_sink_fsm_79_init;
    end else begin
      case(_mystream_sum_vec15_sink_fsm_79)
        _mystream_sum_vec15_sink_fsm_79_init: begin
          if(_mystream_sink_start && _mystream_sum_vec15_sink_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_sum_vec15_sink_fsm_79 <= _mystream_sum_vec15_sink_fsm_79_1;
          end 
        end
        _mystream_sum_vec15_sink_fsm_79_1: begin
          if(_mystream_stream_oready) begin
            _mystream_sum_vec15_sink_fsm_79 <= _mystream_sum_vec15_sink_fsm_79_2;
          end 
        end
        _mystream_sum_vec15_sink_fsm_79_2: begin
          if((_mystream_sum_vec15_sink_count == 1) && _mystream_stream_oready) begin
            _mystream_sum_vec15_sink_fsm_79 <= _mystream_sum_vec15_sink_fsm_79_init;
          end 
          if(_mystream_sink_stop && _mystream_stream_oready) begin
            _mystream_sum_vec15_sink_fsm_79 <= _mystream_sum_vec15_sink_fsm_79_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_sum_vec16_sink_fsm_80_1 = 1;
  localparam _mystream_sum_vec16_sink_fsm_80_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_sum_vec16_sink_fsm_80 <= _mystream_sum_vec16_sink_fsm_80_init;
    end else begin
      case(_mystream_sum_vec16_sink_fsm_80)
        _mystream_sum_vec16_sink_fsm_80_init: begin
          if(_mystream_sink_start && _mystream_sum_vec16_sink_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_sum_vec16_sink_fsm_80 <= _mystream_sum_vec16_sink_fsm_80_1;
          end 
        end
        _mystream_sum_vec16_sink_fsm_80_1: begin
          if(_mystream_stream_oready) begin
            _mystream_sum_vec16_sink_fsm_80 <= _mystream_sum_vec16_sink_fsm_80_2;
          end 
        end
        _mystream_sum_vec16_sink_fsm_80_2: begin
          if((_mystream_sum_vec16_sink_count == 1) && _mystream_stream_oready) begin
            _mystream_sum_vec16_sink_fsm_80 <= _mystream_sum_vec16_sink_fsm_80_init;
          end 
          if(_mystream_sink_stop && _mystream_stream_oready) begin
            _mystream_sum_vec16_sink_fsm_80 <= _mystream_sum_vec16_sink_fsm_80_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_sum_vec17_sink_fsm_81_1 = 1;
  localparam _mystream_sum_vec17_sink_fsm_81_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_sum_vec17_sink_fsm_81 <= _mystream_sum_vec17_sink_fsm_81_init;
    end else begin
      case(_mystream_sum_vec17_sink_fsm_81)
        _mystream_sum_vec17_sink_fsm_81_init: begin
          if(_mystream_sink_start && _mystream_sum_vec17_sink_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_sum_vec17_sink_fsm_81 <= _mystream_sum_vec17_sink_fsm_81_1;
          end 
        end
        _mystream_sum_vec17_sink_fsm_81_1: begin
          if(_mystream_stream_oready) begin
            _mystream_sum_vec17_sink_fsm_81 <= _mystream_sum_vec17_sink_fsm_81_2;
          end 
        end
        _mystream_sum_vec17_sink_fsm_81_2: begin
          if((_mystream_sum_vec17_sink_count == 1) && _mystream_stream_oready) begin
            _mystream_sum_vec17_sink_fsm_81 <= _mystream_sum_vec17_sink_fsm_81_init;
          end 
          if(_mystream_sink_stop && _mystream_stream_oready) begin
            _mystream_sum_vec17_sink_fsm_81 <= _mystream_sum_vec17_sink_fsm_81_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_sum_vec18_sink_fsm_82_1 = 1;
  localparam _mystream_sum_vec18_sink_fsm_82_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_sum_vec18_sink_fsm_82 <= _mystream_sum_vec18_sink_fsm_82_init;
    end else begin
      case(_mystream_sum_vec18_sink_fsm_82)
        _mystream_sum_vec18_sink_fsm_82_init: begin
          if(_mystream_sink_start && _mystream_sum_vec18_sink_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_sum_vec18_sink_fsm_82 <= _mystream_sum_vec18_sink_fsm_82_1;
          end 
        end
        _mystream_sum_vec18_sink_fsm_82_1: begin
          if(_mystream_stream_oready) begin
            _mystream_sum_vec18_sink_fsm_82 <= _mystream_sum_vec18_sink_fsm_82_2;
          end 
        end
        _mystream_sum_vec18_sink_fsm_82_2: begin
          if((_mystream_sum_vec18_sink_count == 1) && _mystream_stream_oready) begin
            _mystream_sum_vec18_sink_fsm_82 <= _mystream_sum_vec18_sink_fsm_82_init;
          end 
          if(_mystream_sink_stop && _mystream_stream_oready) begin
            _mystream_sum_vec18_sink_fsm_82 <= _mystream_sum_vec18_sink_fsm_82_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_sum_vec19_sink_fsm_83_1 = 1;
  localparam _mystream_sum_vec19_sink_fsm_83_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_sum_vec19_sink_fsm_83 <= _mystream_sum_vec19_sink_fsm_83_init;
    end else begin
      case(_mystream_sum_vec19_sink_fsm_83)
        _mystream_sum_vec19_sink_fsm_83_init: begin
          if(_mystream_sink_start && _mystream_sum_vec19_sink_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_sum_vec19_sink_fsm_83 <= _mystream_sum_vec19_sink_fsm_83_1;
          end 
        end
        _mystream_sum_vec19_sink_fsm_83_1: begin
          if(_mystream_stream_oready) begin
            _mystream_sum_vec19_sink_fsm_83 <= _mystream_sum_vec19_sink_fsm_83_2;
          end 
        end
        _mystream_sum_vec19_sink_fsm_83_2: begin
          if((_mystream_sum_vec19_sink_count == 1) && _mystream_stream_oready) begin
            _mystream_sum_vec19_sink_fsm_83 <= _mystream_sum_vec19_sink_fsm_83_init;
          end 
          if(_mystream_sink_stop && _mystream_stream_oready) begin
            _mystream_sum_vec19_sink_fsm_83 <= _mystream_sum_vec19_sink_fsm_83_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_sum_vec20_sink_fsm_84_1 = 1;
  localparam _mystream_sum_vec20_sink_fsm_84_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_sum_vec20_sink_fsm_84 <= _mystream_sum_vec20_sink_fsm_84_init;
    end else begin
      case(_mystream_sum_vec20_sink_fsm_84)
        _mystream_sum_vec20_sink_fsm_84_init: begin
          if(_mystream_sink_start && _mystream_sum_vec20_sink_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_sum_vec20_sink_fsm_84 <= _mystream_sum_vec20_sink_fsm_84_1;
          end 
        end
        _mystream_sum_vec20_sink_fsm_84_1: begin
          if(_mystream_stream_oready) begin
            _mystream_sum_vec20_sink_fsm_84 <= _mystream_sum_vec20_sink_fsm_84_2;
          end 
        end
        _mystream_sum_vec20_sink_fsm_84_2: begin
          if((_mystream_sum_vec20_sink_count == 1) && _mystream_stream_oready) begin
            _mystream_sum_vec20_sink_fsm_84 <= _mystream_sum_vec20_sink_fsm_84_init;
          end 
          if(_mystream_sink_stop && _mystream_stream_oready) begin
            _mystream_sum_vec20_sink_fsm_84 <= _mystream_sum_vec20_sink_fsm_84_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_sum_vec21_sink_fsm_85_1 = 1;
  localparam _mystream_sum_vec21_sink_fsm_85_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_sum_vec21_sink_fsm_85 <= _mystream_sum_vec21_sink_fsm_85_init;
    end else begin
      case(_mystream_sum_vec21_sink_fsm_85)
        _mystream_sum_vec21_sink_fsm_85_init: begin
          if(_mystream_sink_start && _mystream_sum_vec21_sink_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_sum_vec21_sink_fsm_85 <= _mystream_sum_vec21_sink_fsm_85_1;
          end 
        end
        _mystream_sum_vec21_sink_fsm_85_1: begin
          if(_mystream_stream_oready) begin
            _mystream_sum_vec21_sink_fsm_85 <= _mystream_sum_vec21_sink_fsm_85_2;
          end 
        end
        _mystream_sum_vec21_sink_fsm_85_2: begin
          if((_mystream_sum_vec21_sink_count == 1) && _mystream_stream_oready) begin
            _mystream_sum_vec21_sink_fsm_85 <= _mystream_sum_vec21_sink_fsm_85_init;
          end 
          if(_mystream_sink_stop && _mystream_stream_oready) begin
            _mystream_sum_vec21_sink_fsm_85 <= _mystream_sum_vec21_sink_fsm_85_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_sum_vec22_sink_fsm_86_1 = 1;
  localparam _mystream_sum_vec22_sink_fsm_86_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_sum_vec22_sink_fsm_86 <= _mystream_sum_vec22_sink_fsm_86_init;
    end else begin
      case(_mystream_sum_vec22_sink_fsm_86)
        _mystream_sum_vec22_sink_fsm_86_init: begin
          if(_mystream_sink_start && _mystream_sum_vec22_sink_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_sum_vec22_sink_fsm_86 <= _mystream_sum_vec22_sink_fsm_86_1;
          end 
        end
        _mystream_sum_vec22_sink_fsm_86_1: begin
          if(_mystream_stream_oready) begin
            _mystream_sum_vec22_sink_fsm_86 <= _mystream_sum_vec22_sink_fsm_86_2;
          end 
        end
        _mystream_sum_vec22_sink_fsm_86_2: begin
          if((_mystream_sum_vec22_sink_count == 1) && _mystream_stream_oready) begin
            _mystream_sum_vec22_sink_fsm_86 <= _mystream_sum_vec22_sink_fsm_86_init;
          end 
          if(_mystream_sink_stop && _mystream_stream_oready) begin
            _mystream_sum_vec22_sink_fsm_86 <= _mystream_sum_vec22_sink_fsm_86_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_sum_vec23_sink_fsm_87_1 = 1;
  localparam _mystream_sum_vec23_sink_fsm_87_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_sum_vec23_sink_fsm_87 <= _mystream_sum_vec23_sink_fsm_87_init;
    end else begin
      case(_mystream_sum_vec23_sink_fsm_87)
        _mystream_sum_vec23_sink_fsm_87_init: begin
          if(_mystream_sink_start && _mystream_sum_vec23_sink_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_sum_vec23_sink_fsm_87 <= _mystream_sum_vec23_sink_fsm_87_1;
          end 
        end
        _mystream_sum_vec23_sink_fsm_87_1: begin
          if(_mystream_stream_oready) begin
            _mystream_sum_vec23_sink_fsm_87 <= _mystream_sum_vec23_sink_fsm_87_2;
          end 
        end
        _mystream_sum_vec23_sink_fsm_87_2: begin
          if((_mystream_sum_vec23_sink_count == 1) && _mystream_stream_oready) begin
            _mystream_sum_vec23_sink_fsm_87 <= _mystream_sum_vec23_sink_fsm_87_init;
          end 
          if(_mystream_sink_stop && _mystream_stream_oready) begin
            _mystream_sum_vec23_sink_fsm_87 <= _mystream_sum_vec23_sink_fsm_87_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_sum_vec24_sink_fsm_88_1 = 1;
  localparam _mystream_sum_vec24_sink_fsm_88_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_sum_vec24_sink_fsm_88 <= _mystream_sum_vec24_sink_fsm_88_init;
    end else begin
      case(_mystream_sum_vec24_sink_fsm_88)
        _mystream_sum_vec24_sink_fsm_88_init: begin
          if(_mystream_sink_start && _mystream_sum_vec24_sink_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_sum_vec24_sink_fsm_88 <= _mystream_sum_vec24_sink_fsm_88_1;
          end 
        end
        _mystream_sum_vec24_sink_fsm_88_1: begin
          if(_mystream_stream_oready) begin
            _mystream_sum_vec24_sink_fsm_88 <= _mystream_sum_vec24_sink_fsm_88_2;
          end 
        end
        _mystream_sum_vec24_sink_fsm_88_2: begin
          if((_mystream_sum_vec24_sink_count == 1) && _mystream_stream_oready) begin
            _mystream_sum_vec24_sink_fsm_88 <= _mystream_sum_vec24_sink_fsm_88_init;
          end 
          if(_mystream_sink_stop && _mystream_stream_oready) begin
            _mystream_sum_vec24_sink_fsm_88 <= _mystream_sum_vec24_sink_fsm_88_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_sum_vec25_sink_fsm_89_1 = 1;
  localparam _mystream_sum_vec25_sink_fsm_89_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_sum_vec25_sink_fsm_89 <= _mystream_sum_vec25_sink_fsm_89_init;
    end else begin
      case(_mystream_sum_vec25_sink_fsm_89)
        _mystream_sum_vec25_sink_fsm_89_init: begin
          if(_mystream_sink_start && _mystream_sum_vec25_sink_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_sum_vec25_sink_fsm_89 <= _mystream_sum_vec25_sink_fsm_89_1;
          end 
        end
        _mystream_sum_vec25_sink_fsm_89_1: begin
          if(_mystream_stream_oready) begin
            _mystream_sum_vec25_sink_fsm_89 <= _mystream_sum_vec25_sink_fsm_89_2;
          end 
        end
        _mystream_sum_vec25_sink_fsm_89_2: begin
          if((_mystream_sum_vec25_sink_count == 1) && _mystream_stream_oready) begin
            _mystream_sum_vec25_sink_fsm_89 <= _mystream_sum_vec25_sink_fsm_89_init;
          end 
          if(_mystream_sink_stop && _mystream_stream_oready) begin
            _mystream_sum_vec25_sink_fsm_89 <= _mystream_sum_vec25_sink_fsm_89_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_sum_vec26_sink_fsm_90_1 = 1;
  localparam _mystream_sum_vec26_sink_fsm_90_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_sum_vec26_sink_fsm_90 <= _mystream_sum_vec26_sink_fsm_90_init;
    end else begin
      case(_mystream_sum_vec26_sink_fsm_90)
        _mystream_sum_vec26_sink_fsm_90_init: begin
          if(_mystream_sink_start && _mystream_sum_vec26_sink_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_sum_vec26_sink_fsm_90 <= _mystream_sum_vec26_sink_fsm_90_1;
          end 
        end
        _mystream_sum_vec26_sink_fsm_90_1: begin
          if(_mystream_stream_oready) begin
            _mystream_sum_vec26_sink_fsm_90 <= _mystream_sum_vec26_sink_fsm_90_2;
          end 
        end
        _mystream_sum_vec26_sink_fsm_90_2: begin
          if((_mystream_sum_vec26_sink_count == 1) && _mystream_stream_oready) begin
            _mystream_sum_vec26_sink_fsm_90 <= _mystream_sum_vec26_sink_fsm_90_init;
          end 
          if(_mystream_sink_stop && _mystream_stream_oready) begin
            _mystream_sum_vec26_sink_fsm_90 <= _mystream_sum_vec26_sink_fsm_90_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_sum_vec27_sink_fsm_91_1 = 1;
  localparam _mystream_sum_vec27_sink_fsm_91_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_sum_vec27_sink_fsm_91 <= _mystream_sum_vec27_sink_fsm_91_init;
    end else begin
      case(_mystream_sum_vec27_sink_fsm_91)
        _mystream_sum_vec27_sink_fsm_91_init: begin
          if(_mystream_sink_start && _mystream_sum_vec27_sink_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_sum_vec27_sink_fsm_91 <= _mystream_sum_vec27_sink_fsm_91_1;
          end 
        end
        _mystream_sum_vec27_sink_fsm_91_1: begin
          if(_mystream_stream_oready) begin
            _mystream_sum_vec27_sink_fsm_91 <= _mystream_sum_vec27_sink_fsm_91_2;
          end 
        end
        _mystream_sum_vec27_sink_fsm_91_2: begin
          if((_mystream_sum_vec27_sink_count == 1) && _mystream_stream_oready) begin
            _mystream_sum_vec27_sink_fsm_91 <= _mystream_sum_vec27_sink_fsm_91_init;
          end 
          if(_mystream_sink_stop && _mystream_stream_oready) begin
            _mystream_sum_vec27_sink_fsm_91 <= _mystream_sum_vec27_sink_fsm_91_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_sum_vec28_sink_fsm_92_1 = 1;
  localparam _mystream_sum_vec28_sink_fsm_92_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_sum_vec28_sink_fsm_92 <= _mystream_sum_vec28_sink_fsm_92_init;
    end else begin
      case(_mystream_sum_vec28_sink_fsm_92)
        _mystream_sum_vec28_sink_fsm_92_init: begin
          if(_mystream_sink_start && _mystream_sum_vec28_sink_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_sum_vec28_sink_fsm_92 <= _mystream_sum_vec28_sink_fsm_92_1;
          end 
        end
        _mystream_sum_vec28_sink_fsm_92_1: begin
          if(_mystream_stream_oready) begin
            _mystream_sum_vec28_sink_fsm_92 <= _mystream_sum_vec28_sink_fsm_92_2;
          end 
        end
        _mystream_sum_vec28_sink_fsm_92_2: begin
          if((_mystream_sum_vec28_sink_count == 1) && _mystream_stream_oready) begin
            _mystream_sum_vec28_sink_fsm_92 <= _mystream_sum_vec28_sink_fsm_92_init;
          end 
          if(_mystream_sink_stop && _mystream_stream_oready) begin
            _mystream_sum_vec28_sink_fsm_92 <= _mystream_sum_vec28_sink_fsm_92_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_sum_vec29_sink_fsm_93_1 = 1;
  localparam _mystream_sum_vec29_sink_fsm_93_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_sum_vec29_sink_fsm_93 <= _mystream_sum_vec29_sink_fsm_93_init;
    end else begin
      case(_mystream_sum_vec29_sink_fsm_93)
        _mystream_sum_vec29_sink_fsm_93_init: begin
          if(_mystream_sink_start && _mystream_sum_vec29_sink_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_sum_vec29_sink_fsm_93 <= _mystream_sum_vec29_sink_fsm_93_1;
          end 
        end
        _mystream_sum_vec29_sink_fsm_93_1: begin
          if(_mystream_stream_oready) begin
            _mystream_sum_vec29_sink_fsm_93 <= _mystream_sum_vec29_sink_fsm_93_2;
          end 
        end
        _mystream_sum_vec29_sink_fsm_93_2: begin
          if((_mystream_sum_vec29_sink_count == 1) && _mystream_stream_oready) begin
            _mystream_sum_vec29_sink_fsm_93 <= _mystream_sum_vec29_sink_fsm_93_init;
          end 
          if(_mystream_sink_stop && _mystream_stream_oready) begin
            _mystream_sum_vec29_sink_fsm_93 <= _mystream_sum_vec29_sink_fsm_93_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_sum_vec30_sink_fsm_94_1 = 1;
  localparam _mystream_sum_vec30_sink_fsm_94_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_sum_vec30_sink_fsm_94 <= _mystream_sum_vec30_sink_fsm_94_init;
    end else begin
      case(_mystream_sum_vec30_sink_fsm_94)
        _mystream_sum_vec30_sink_fsm_94_init: begin
          if(_mystream_sink_start && _mystream_sum_vec30_sink_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_sum_vec30_sink_fsm_94 <= _mystream_sum_vec30_sink_fsm_94_1;
          end 
        end
        _mystream_sum_vec30_sink_fsm_94_1: begin
          if(_mystream_stream_oready) begin
            _mystream_sum_vec30_sink_fsm_94 <= _mystream_sum_vec30_sink_fsm_94_2;
          end 
        end
        _mystream_sum_vec30_sink_fsm_94_2: begin
          if((_mystream_sum_vec30_sink_count == 1) && _mystream_stream_oready) begin
            _mystream_sum_vec30_sink_fsm_94 <= _mystream_sum_vec30_sink_fsm_94_init;
          end 
          if(_mystream_sink_stop && _mystream_stream_oready) begin
            _mystream_sum_vec30_sink_fsm_94 <= _mystream_sum_vec30_sink_fsm_94_init;
          end 
        end
      endcase
    end
  end

  localparam _mystream_sum_vec31_sink_fsm_95_1 = 1;
  localparam _mystream_sum_vec31_sink_fsm_95_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _mystream_sum_vec31_sink_fsm_95 <= _mystream_sum_vec31_sink_fsm_95_init;
    end else begin
      case(_mystream_sum_vec31_sink_fsm_95)
        _mystream_sum_vec31_sink_fsm_95_init: begin
          if(_mystream_sink_start && _mystream_sum_vec31_sink_mode & 5'b1 && _mystream_stream_oready) begin
            _mystream_sum_vec31_sink_fsm_95 <= _mystream_sum_vec31_sink_fsm_95_1;
          end 
        end
        _mystream_sum_vec31_sink_fsm_95_1: begin
          if(_mystream_stream_oready) begin
            _mystream_sum_vec31_sink_fsm_95 <= _mystream_sum_vec31_sink_fsm_95_2;
          end 
        end
        _mystream_sum_vec31_sink_fsm_95_2: begin
          if((_mystream_sum_vec31_sink_count == 1) && _mystream_stream_oready) begin
            _mystream_sum_vec31_sink_fsm_95 <= _mystream_sum_vec31_sink_fsm_95_init;
          end 
          if(_mystream_sink_stop && _mystream_stream_oready) begin
            _mystream_sum_vec31_sink_fsm_95 <= _mystream_sum_vec31_sink_fsm_95_init;
          end 
        end
      endcase
    end
  end

  localparam _myaxi_read_data_fsm_1 = 1;
  localparam _myaxi_read_data_fsm_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _myaxi_read_data_fsm <= _myaxi_read_data_fsm_init;
    end else begin
      case(_myaxi_read_data_fsm)
        _myaxi_read_data_fsm_init: begin
          if(_myaxi_read_data_idle && !_myaxi_read_req_fifo_empty && (_myaxi_read_op_sel_fifo == 3)) begin
            _myaxi_read_data_fsm <= _myaxi_read_data_fsm_1;
          end 
          if(_myaxi_read_data_idle && !_myaxi_read_req_fifo_empty && (_myaxi_read_op_sel_fifo == 4)) begin
            _myaxi_read_data_fsm <= _myaxi_read_data_fsm_1;
          end 
        end
        _myaxi_read_data_fsm_1: begin
          _myaxi_read_data_fsm <= _myaxi_read_data_fsm_2;
          _myaxi_read_data_fsm <= _myaxi_read_data_fsm_2;
        end
        _myaxi_read_data_fsm_2: begin
          if(myaxi_rvalid && (_myaxi_read_local_size_buf <= 1)) begin
            _myaxi_read_data_fsm <= _myaxi_read_data_fsm_init;
          end 
          if(myaxi_rvalid && (_myaxi_read_local_size_buf <= 1)) begin
            _myaxi_read_data_fsm <= _myaxi_read_data_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_2_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_2 <= write_burst_fsm_2_init;
      write_burst_addr_1087 <= 0;
      write_burst_stride_1088 <= 0;
      write_burst_length_1089 <= 0;
      write_burst_done_1090 <= 0;
    end else begin
      case(write_burst_fsm_2)
        write_burst_fsm_2_init: begin
          write_burst_addr_1087 <= _myaxi_read_local_addr_buf;
          write_burst_stride_1088 <= _myaxi_read_local_stride_buf;
          write_burst_length_1089 <= _myaxi_read_local_size_buf;
          write_burst_done_1090 <= 0;
          if((_myaxi_read_data_fsm == 1) && (_myaxi_read_op_sel_buf == 3) && (_myaxi_read_local_size_buf > 0)) begin
            write_burst_fsm_2 <= write_burst_fsm_2_1;
          end 
        end
        write_burst_fsm_2_1: begin
          if(myaxi_rvalid) begin
            write_burst_addr_1087 <= write_burst_addr_1087 + write_burst_stride_1088;
            write_burst_length_1089 <= write_burst_length_1089 - 1;
            write_burst_done_1090 <= 0;
          end 
          if(myaxi_rvalid && (write_burst_length_1089 <= 1)) begin
            write_burst_done_1090 <= 1;
          end 
          if(myaxi_rvalid && 0) begin
            write_burst_done_1090 <= 1;
          end 
          if(myaxi_rvalid && (write_burst_length_1089 <= 1)) begin
            write_burst_fsm_2 <= write_burst_fsm_2_init;
          end 
          if(myaxi_rvalid && 0) begin
            write_burst_fsm_2 <= write_burst_fsm_2_init;
          end 
          if(0) begin
            write_burst_fsm_2 <= write_burst_fsm_2_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_fsm_3_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_fsm_3 <= write_burst_fsm_3_init;
      write_burst_addr_1093 <= 0;
      write_burst_stride_1094 <= 0;
      write_burst_length_1095 <= 0;
      write_burst_done_1096 <= 0;
    end else begin
      case(write_burst_fsm_3)
        write_burst_fsm_3_init: begin
          write_burst_addr_1093 <= _myaxi_read_local_addr_buf;
          write_burst_stride_1094 <= _myaxi_read_local_stride_buf;
          write_burst_length_1095 <= _myaxi_read_local_size_buf;
          write_burst_done_1096 <= 0;
          if((_myaxi_read_data_fsm == 1) && (_myaxi_read_op_sel_buf == 4) && (_myaxi_read_local_size_buf > 0)) begin
            write_burst_fsm_3 <= write_burst_fsm_3_1;
          end 
        end
        write_burst_fsm_3_1: begin
          if(myaxi_rvalid) begin
            write_burst_addr_1093 <= write_burst_addr_1093 + write_burst_stride_1094;
            write_burst_length_1095 <= write_burst_length_1095 - 1;
            write_burst_done_1096 <= 0;
          end 
          if(myaxi_rvalid && (write_burst_length_1095 <= 1)) begin
            write_burst_done_1096 <= 1;
          end 
          if(myaxi_rvalid && 0) begin
            write_burst_done_1096 <= 1;
          end 
          if(myaxi_rvalid && (write_burst_length_1095 <= 1)) begin
            write_burst_fsm_3 <= write_burst_fsm_3_init;
          end 
          if(myaxi_rvalid && 0) begin
            write_burst_fsm_3 <= write_burst_fsm_3_init;
          end 
          if(0) begin
            write_burst_fsm_3 <= write_burst_fsm_3_init;
          end 
        end
      endcase
    end
  end

  localparam _myaxi_write_req_fsm_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      _myaxi_write_req_fsm <= _myaxi_write_req_fsm_init;
      _myaxi_write_cont <= 0;
    end else begin
      case(_myaxi_write_req_fsm)
        _myaxi_write_req_fsm_init: begin
          if((_myaxi_write_req_fsm == 0) && (_myaxi_write_start || _myaxi_write_cont) && !_myaxi_write_req_fifo_almost_full) begin
            _myaxi_write_req_fsm <= _myaxi_write_req_fsm_1;
          end 
        end
        _myaxi_write_req_fsm_1: begin
          if((_myaxi_write_req_fsm == 1) && !_myaxi_write_req_fifo_almost_full && (myaxi_awready || !myaxi_awvalid) && (outstanding_wcount_0 < 6)) begin
            _myaxi_write_cont <= 1;
          end 
          if((_myaxi_write_req_fsm == 1) && !_myaxi_write_req_fifo_almost_full && (myaxi_awready || !myaxi_awvalid) && (outstanding_wcount_0 < 6) && (_myaxi_write_global_size == 0)) begin
            _myaxi_write_cont <= 0;
          end 
          if((_myaxi_write_req_fsm == 1) && !_myaxi_write_req_fifo_almost_full && (myaxi_awready || !myaxi_awvalid) && (outstanding_wcount_0 < 6)) begin
            _myaxi_write_req_fsm <= _myaxi_write_req_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam _myaxi_write_data_fsm_1 = 1;
  localparam _myaxi_write_data_fsm_2 = 2;

  always @(posedge CLK) begin
    if(RST) begin
      _myaxi_write_data_fsm <= _myaxi_write_data_fsm_init;
    end else begin
      case(_myaxi_write_data_fsm)
        _myaxi_write_data_fsm_init: begin
          if(_myaxi_write_data_idle && !_myaxi_write_req_fifo_empty && (_myaxi_write_op_sel_fifo == 1)) begin
            _myaxi_write_data_fsm <= _myaxi_write_data_fsm_1;
          end 
        end
        _myaxi_write_data_fsm_1: begin
          _myaxi_write_data_fsm <= _myaxi_write_data_fsm_2;
        end
        _myaxi_write_data_fsm_2: begin
          if((_myaxi_write_op_sel_buf == 1) && read_burst_rvalid_1136 && ((myaxi_wready || !myaxi_wvalid) && (_myaxi_write_size_buf > 0)) && read_burst_rlast_1137) begin
            _myaxi_write_data_fsm <= _myaxi_write_data_fsm_init;
          end 
        end
      endcase
    end
  end

  localparam read_burst_fsm_4_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      read_burst_fsm_4 <= read_burst_fsm_4_init;
      read_burst_addr_1133 <= 0;
      read_burst_stride_1134 <= 0;
      read_burst_length_1135 <= 0;
      read_burst_rvalid_1136 <= 0;
      read_burst_rlast_1137 <= 0;
    end else begin
      case(read_burst_fsm_4)
        read_burst_fsm_4_init: begin
          read_burst_addr_1133 <= _myaxi_write_local_addr_buf;
          read_burst_stride_1134 <= _myaxi_write_local_stride_buf;
          read_burst_length_1135 <= _myaxi_write_size_buf;
          read_burst_rvalid_1136 <= 0;
          read_burst_rlast_1137 <= 0;
          if((_myaxi_write_data_fsm == 1) && (_myaxi_write_op_sel_buf == 1) && (_myaxi_write_size_buf > 0)) begin
            read_burst_fsm_4 <= read_burst_fsm_4_1;
          end 
        end
        read_burst_fsm_4_1: begin
          if((myaxi_wready || !myaxi_wvalid) && (_myaxi_write_size_buf > 0) && (read_burst_length_1135 > 0)) begin
            read_burst_addr_1133 <= read_burst_addr_1133 + read_burst_stride_1134;
            read_burst_length_1135 <= read_burst_length_1135 - 1;
            read_burst_rvalid_1136 <= 1;
          end 
          if((myaxi_wready || !myaxi_wvalid) && (_myaxi_write_size_buf > 0) && (read_burst_length_1135 <= 1)) begin
            read_burst_rlast_1137 <= 1;
          end 
          if(read_burst_rlast_1137 && read_burst_rvalid_1136 && ((myaxi_wready || !myaxi_wvalid) && (_myaxi_write_size_buf > 0))) begin
            read_burst_rvalid_1136 <= 0;
            read_burst_rlast_1137 <= 0;
          end 
          if(0) begin
            read_burst_rvalid_1136 <= 0;
            read_burst_rlast_1137 <= 0;
          end 
          if(read_burst_rlast_1137 && read_burst_rvalid_1136 && ((myaxi_wready || !myaxi_wvalid) && (_myaxi_write_size_buf > 0))) begin
            read_burst_fsm_4 <= read_burst_fsm_4_init;
          end 
          if(0) begin
            read_burst_fsm_4 <= read_burst_fsm_4_init;
          end 
        end
      endcase
    end
  end

  localparam write_burst_packed_fsm_5_1 = 1;

  always @(posedge CLK) begin
    if(RST) begin
      write_burst_packed_fsm_5 <= write_burst_packed_fsm_5_init;
      write_burst_packed_addr_1149 <= 0;
      write_burst_packed_stride_1150 <= 0;
      write_burst_packed_length_1151 <= 0;
      write_burst_packed_done_1152 <= 0;
    end else begin
      case(write_burst_packed_fsm_5)
        write_burst_packed_fsm_5_init: begin
          write_burst_packed_addr_1149 <= _myaxi_read_local_addr_buf;
          write_burst_packed_stride_1150 <= _myaxi_read_local_stride_buf;
          write_burst_packed_length_1151 <= _myaxi_read_local_size_buf;
          write_burst_packed_done_1152 <= 0;
          if((_myaxi_read_data_narrow_fsm == 1) && (_myaxi_read_op_sel_buf == 5) && (_myaxi_read_local_size_buf > 0)) begin
            write_burst_packed_fsm_5 <= write_burst_packed_fsm_5_1;
          end 
        end
        write_burst_packed_fsm_5_1: begin
          if(_myaxi_read_narrow_wvalid_1147) begin
            write_burst_packed_addr_1149 <= write_burst_packed_addr_1149 + write_burst_packed_stride_1150;
            write_burst_packed_length_1151 <= write_burst_packed_length_1151 - 1;
            write_burst_packed_done_1152 <= 0;
          end 
          if(_myaxi_read_narrow_wvalid_1147 && (write_burst_packed_length_1151 <= 1)) begin
            write_burst_packed_done_1152 <= 1;
          end 
          if(_myaxi_read_narrow_wvalid_1147 && 0) begin
            write_burst_packed_done_1152 <= 1;
          end 
          if(_myaxi_read_narrow_wvalid_1147 && (write_burst_packed_length_1151 <= 1)) begin
            write_burst_packed_fsm_5 <= write_burst_packed_fsm_5_init;
          end 
          if(_myaxi_read_narrow_wvalid_1147 && 0) begin
            write_burst_packed_fsm_5 <= write_burst_packed_fsm_5_init;
          end 
          if(0) begin
            write_burst_packed_fsm_5 <= write_burst_packed_fsm_5_init;
          end 
        end
      endcase
    end
  end


  always @(posedge CLK) begin
    if(RST) begin
      _tmp_1218 <= 0;
      _tmp_1287 <= 0;
    end else begin
      if(th_comp == 114) begin
        _tmp_1218 <= read_rtl_bank_1217;
      end 
      if(th_comp == 116) begin
        _tmp_1287 <= read_rtl_bank_1286;
      end 
    end
  end


endmodule



module _myaxi_read_req_fifo
(
  input CLK,
  input RST,
  input _myaxi_read_req_fifo_enq,
  input [137-1:0] _myaxi_read_req_fifo_wdata,
  output _myaxi_read_req_fifo_full,
  output _myaxi_read_req_fifo_almost_full,
  input _myaxi_read_req_fifo_deq,
  output [137-1:0] _myaxi_read_req_fifo_rdata,
  output _myaxi_read_req_fifo_empty,
  output _myaxi_read_req_fifo_almost_empty
);

  reg [137-1:0] mem [0:8-1];
  reg [3-1:0] head;
  reg [3-1:0] tail;
  wire is_empty;
  wire is_almost_empty;
  wire is_full;
  wire is_almost_full;
  assign is_empty = head == tail;
  assign is_almost_empty = head == (tail + 1 & 7);
  assign is_full = (head + 1 & 7) == tail;
  assign is_almost_full = (head + 2 & 7) == tail;
  wire [137-1:0] rdata;
  assign _myaxi_read_req_fifo_full = is_full;
  assign _myaxi_read_req_fifo_almost_full = is_almost_full || is_full;
  assign _myaxi_read_req_fifo_empty = is_empty;
  assign _myaxi_read_req_fifo_almost_empty = is_almost_empty || is_empty;
  assign rdata = mem[tail];
  assign _myaxi_read_req_fifo_rdata = rdata;

  always @(posedge CLK) begin
    if(RST) begin
      head <= 0;
      tail <= 0;
    end else begin
      if(_myaxi_read_req_fifo_enq && !is_full) begin
        mem[head] <= _myaxi_read_req_fifo_wdata;
        head <= head + 1;
      end 
      if(_myaxi_read_req_fifo_deq && !is_empty) begin
        tail <= tail + 1;
      end 
    end
  end


endmodule



module _myaxi_write_req_fifo
(
  input CLK,
  input RST,
  input _myaxi_write_req_fifo_enq,
  input [137-1:0] _myaxi_write_req_fifo_wdata,
  output _myaxi_write_req_fifo_full,
  output _myaxi_write_req_fifo_almost_full,
  input _myaxi_write_req_fifo_deq,
  output [137-1:0] _myaxi_write_req_fifo_rdata,
  output _myaxi_write_req_fifo_empty,
  output _myaxi_write_req_fifo_almost_empty
);

  reg [137-1:0] mem [0:8-1];
  reg [3-1:0] head;
  reg [3-1:0] tail;
  wire is_empty;
  wire is_almost_empty;
  wire is_full;
  wire is_almost_full;
  assign is_empty = head == tail;
  assign is_almost_empty = head == (tail + 1 & 7);
  assign is_full = (head + 1 & 7) == tail;
  assign is_almost_full = (head + 2 & 7) == tail;
  wire [137-1:0] rdata;
  assign _myaxi_write_req_fifo_full = is_full;
  assign _myaxi_write_req_fifo_almost_full = is_almost_full || is_full;
  assign _myaxi_write_req_fifo_empty = is_empty;
  assign _myaxi_write_req_fifo_almost_empty = is_almost_empty || is_empty;
  assign rdata = mem[tail];
  assign _myaxi_write_req_fifo_rdata = rdata;

  always @(posedge CLK) begin
    if(RST) begin
      head <= 0;
      tail <= 0;
    end else begin
      if(_myaxi_write_req_fifo_enq && !is_full) begin
        mem[head] <= _myaxi_write_req_fifo_wdata;
        head <= head + 1;
      end 
      if(_myaxi_write_req_fifo_deq && !is_empty) begin
        tail <= tail + 1;
      end 
    end
  end


endmodule



module ram_a_0
(
  input CLK,
  input [20-1:0] ram_a_0_0_addr,
  output [32-1:0] ram_a_0_0_rdata,
  input [32-1:0] ram_a_0_0_wdata,
  input ram_a_0_0_wenable,
  input ram_a_0_0_enable
);

  reg [32-1:0] ram_a_0_0_rdata_out;
  assign ram_a_0_0_rdata = ram_a_0_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_a_0_0_enable) begin
      if(ram_a_0_0_wenable) begin
        mem[ram_a_0_0_addr] <= ram_a_0_0_wdata;
        ram_a_0_0_rdata_out <= ram_a_0_0_wdata;
      end else begin
        ram_a_0_0_rdata_out <= mem[ram_a_0_0_addr];
      end
    end 
  end


endmodule



module ram_a_1
(
  input CLK,
  input [20-1:0] ram_a_1_0_addr,
  output [32-1:0] ram_a_1_0_rdata,
  input [32-1:0] ram_a_1_0_wdata,
  input ram_a_1_0_wenable,
  input ram_a_1_0_enable
);

  reg [32-1:0] ram_a_1_0_rdata_out;
  assign ram_a_1_0_rdata = ram_a_1_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_a_1_0_enable) begin
      if(ram_a_1_0_wenable) begin
        mem[ram_a_1_0_addr] <= ram_a_1_0_wdata;
        ram_a_1_0_rdata_out <= ram_a_1_0_wdata;
      end else begin
        ram_a_1_0_rdata_out <= mem[ram_a_1_0_addr];
      end
    end 
  end


endmodule



module ram_a_2
(
  input CLK,
  input [20-1:0] ram_a_2_0_addr,
  output [32-1:0] ram_a_2_0_rdata,
  input [32-1:0] ram_a_2_0_wdata,
  input ram_a_2_0_wenable,
  input ram_a_2_0_enable
);

  reg [32-1:0] ram_a_2_0_rdata_out;
  assign ram_a_2_0_rdata = ram_a_2_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_a_2_0_enable) begin
      if(ram_a_2_0_wenable) begin
        mem[ram_a_2_0_addr] <= ram_a_2_0_wdata;
        ram_a_2_0_rdata_out <= ram_a_2_0_wdata;
      end else begin
        ram_a_2_0_rdata_out <= mem[ram_a_2_0_addr];
      end
    end 
  end


endmodule



module ram_a_3
(
  input CLK,
  input [20-1:0] ram_a_3_0_addr,
  output [32-1:0] ram_a_3_0_rdata,
  input [32-1:0] ram_a_3_0_wdata,
  input ram_a_3_0_wenable,
  input ram_a_3_0_enable
);

  reg [32-1:0] ram_a_3_0_rdata_out;
  assign ram_a_3_0_rdata = ram_a_3_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_a_3_0_enable) begin
      if(ram_a_3_0_wenable) begin
        mem[ram_a_3_0_addr] <= ram_a_3_0_wdata;
        ram_a_3_0_rdata_out <= ram_a_3_0_wdata;
      end else begin
        ram_a_3_0_rdata_out <= mem[ram_a_3_0_addr];
      end
    end 
  end


endmodule



module ram_a_4
(
  input CLK,
  input [20-1:0] ram_a_4_0_addr,
  output [32-1:0] ram_a_4_0_rdata,
  input [32-1:0] ram_a_4_0_wdata,
  input ram_a_4_0_wenable,
  input ram_a_4_0_enable
);

  reg [32-1:0] ram_a_4_0_rdata_out;
  assign ram_a_4_0_rdata = ram_a_4_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_a_4_0_enable) begin
      if(ram_a_4_0_wenable) begin
        mem[ram_a_4_0_addr] <= ram_a_4_0_wdata;
        ram_a_4_0_rdata_out <= ram_a_4_0_wdata;
      end else begin
        ram_a_4_0_rdata_out <= mem[ram_a_4_0_addr];
      end
    end 
  end


endmodule



module ram_a_5
(
  input CLK,
  input [20-1:0] ram_a_5_0_addr,
  output [32-1:0] ram_a_5_0_rdata,
  input [32-1:0] ram_a_5_0_wdata,
  input ram_a_5_0_wenable,
  input ram_a_5_0_enable
);

  reg [32-1:0] ram_a_5_0_rdata_out;
  assign ram_a_5_0_rdata = ram_a_5_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_a_5_0_enable) begin
      if(ram_a_5_0_wenable) begin
        mem[ram_a_5_0_addr] <= ram_a_5_0_wdata;
        ram_a_5_0_rdata_out <= ram_a_5_0_wdata;
      end else begin
        ram_a_5_0_rdata_out <= mem[ram_a_5_0_addr];
      end
    end 
  end


endmodule



module ram_a_6
(
  input CLK,
  input [20-1:0] ram_a_6_0_addr,
  output [32-1:0] ram_a_6_0_rdata,
  input [32-1:0] ram_a_6_0_wdata,
  input ram_a_6_0_wenable,
  input ram_a_6_0_enable
);

  reg [32-1:0] ram_a_6_0_rdata_out;
  assign ram_a_6_0_rdata = ram_a_6_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_a_6_0_enable) begin
      if(ram_a_6_0_wenable) begin
        mem[ram_a_6_0_addr] <= ram_a_6_0_wdata;
        ram_a_6_0_rdata_out <= ram_a_6_0_wdata;
      end else begin
        ram_a_6_0_rdata_out <= mem[ram_a_6_0_addr];
      end
    end 
  end


endmodule



module ram_a_7
(
  input CLK,
  input [20-1:0] ram_a_7_0_addr,
  output [32-1:0] ram_a_7_0_rdata,
  input [32-1:0] ram_a_7_0_wdata,
  input ram_a_7_0_wenable,
  input ram_a_7_0_enable
);

  reg [32-1:0] ram_a_7_0_rdata_out;
  assign ram_a_7_0_rdata = ram_a_7_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_a_7_0_enable) begin
      if(ram_a_7_0_wenable) begin
        mem[ram_a_7_0_addr] <= ram_a_7_0_wdata;
        ram_a_7_0_rdata_out <= ram_a_7_0_wdata;
      end else begin
        ram_a_7_0_rdata_out <= mem[ram_a_7_0_addr];
      end
    end 
  end


endmodule



module ram_a_8
(
  input CLK,
  input [20-1:0] ram_a_8_0_addr,
  output [32-1:0] ram_a_8_0_rdata,
  input [32-1:0] ram_a_8_0_wdata,
  input ram_a_8_0_wenable,
  input ram_a_8_0_enable
);

  reg [32-1:0] ram_a_8_0_rdata_out;
  assign ram_a_8_0_rdata = ram_a_8_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_a_8_0_enable) begin
      if(ram_a_8_0_wenable) begin
        mem[ram_a_8_0_addr] <= ram_a_8_0_wdata;
        ram_a_8_0_rdata_out <= ram_a_8_0_wdata;
      end else begin
        ram_a_8_0_rdata_out <= mem[ram_a_8_0_addr];
      end
    end 
  end


endmodule



module ram_a_9
(
  input CLK,
  input [20-1:0] ram_a_9_0_addr,
  output [32-1:0] ram_a_9_0_rdata,
  input [32-1:0] ram_a_9_0_wdata,
  input ram_a_9_0_wenable,
  input ram_a_9_0_enable
);

  reg [32-1:0] ram_a_9_0_rdata_out;
  assign ram_a_9_0_rdata = ram_a_9_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_a_9_0_enable) begin
      if(ram_a_9_0_wenable) begin
        mem[ram_a_9_0_addr] <= ram_a_9_0_wdata;
        ram_a_9_0_rdata_out <= ram_a_9_0_wdata;
      end else begin
        ram_a_9_0_rdata_out <= mem[ram_a_9_0_addr];
      end
    end 
  end


endmodule



module ram_a_10
(
  input CLK,
  input [20-1:0] ram_a_10_0_addr,
  output [32-1:0] ram_a_10_0_rdata,
  input [32-1:0] ram_a_10_0_wdata,
  input ram_a_10_0_wenable,
  input ram_a_10_0_enable
);

  reg [32-1:0] ram_a_10_0_rdata_out;
  assign ram_a_10_0_rdata = ram_a_10_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_a_10_0_enable) begin
      if(ram_a_10_0_wenable) begin
        mem[ram_a_10_0_addr] <= ram_a_10_0_wdata;
        ram_a_10_0_rdata_out <= ram_a_10_0_wdata;
      end else begin
        ram_a_10_0_rdata_out <= mem[ram_a_10_0_addr];
      end
    end 
  end


endmodule



module ram_a_11
(
  input CLK,
  input [20-1:0] ram_a_11_0_addr,
  output [32-1:0] ram_a_11_0_rdata,
  input [32-1:0] ram_a_11_0_wdata,
  input ram_a_11_0_wenable,
  input ram_a_11_0_enable
);

  reg [32-1:0] ram_a_11_0_rdata_out;
  assign ram_a_11_0_rdata = ram_a_11_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_a_11_0_enable) begin
      if(ram_a_11_0_wenable) begin
        mem[ram_a_11_0_addr] <= ram_a_11_0_wdata;
        ram_a_11_0_rdata_out <= ram_a_11_0_wdata;
      end else begin
        ram_a_11_0_rdata_out <= mem[ram_a_11_0_addr];
      end
    end 
  end


endmodule



module ram_a_12
(
  input CLK,
  input [20-1:0] ram_a_12_0_addr,
  output [32-1:0] ram_a_12_0_rdata,
  input [32-1:0] ram_a_12_0_wdata,
  input ram_a_12_0_wenable,
  input ram_a_12_0_enable
);

  reg [32-1:0] ram_a_12_0_rdata_out;
  assign ram_a_12_0_rdata = ram_a_12_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_a_12_0_enable) begin
      if(ram_a_12_0_wenable) begin
        mem[ram_a_12_0_addr] <= ram_a_12_0_wdata;
        ram_a_12_0_rdata_out <= ram_a_12_0_wdata;
      end else begin
        ram_a_12_0_rdata_out <= mem[ram_a_12_0_addr];
      end
    end 
  end


endmodule



module ram_a_13
(
  input CLK,
  input [20-1:0] ram_a_13_0_addr,
  output [32-1:0] ram_a_13_0_rdata,
  input [32-1:0] ram_a_13_0_wdata,
  input ram_a_13_0_wenable,
  input ram_a_13_0_enable
);

  reg [32-1:0] ram_a_13_0_rdata_out;
  assign ram_a_13_0_rdata = ram_a_13_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_a_13_0_enable) begin
      if(ram_a_13_0_wenable) begin
        mem[ram_a_13_0_addr] <= ram_a_13_0_wdata;
        ram_a_13_0_rdata_out <= ram_a_13_0_wdata;
      end else begin
        ram_a_13_0_rdata_out <= mem[ram_a_13_0_addr];
      end
    end 
  end


endmodule



module ram_a_14
(
  input CLK,
  input [20-1:0] ram_a_14_0_addr,
  output [32-1:0] ram_a_14_0_rdata,
  input [32-1:0] ram_a_14_0_wdata,
  input ram_a_14_0_wenable,
  input ram_a_14_0_enable
);

  reg [32-1:0] ram_a_14_0_rdata_out;
  assign ram_a_14_0_rdata = ram_a_14_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_a_14_0_enable) begin
      if(ram_a_14_0_wenable) begin
        mem[ram_a_14_0_addr] <= ram_a_14_0_wdata;
        ram_a_14_0_rdata_out <= ram_a_14_0_wdata;
      end else begin
        ram_a_14_0_rdata_out <= mem[ram_a_14_0_addr];
      end
    end 
  end


endmodule



module ram_a_15
(
  input CLK,
  input [20-1:0] ram_a_15_0_addr,
  output [32-1:0] ram_a_15_0_rdata,
  input [32-1:0] ram_a_15_0_wdata,
  input ram_a_15_0_wenable,
  input ram_a_15_0_enable
);

  reg [32-1:0] ram_a_15_0_rdata_out;
  assign ram_a_15_0_rdata = ram_a_15_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_a_15_0_enable) begin
      if(ram_a_15_0_wenable) begin
        mem[ram_a_15_0_addr] <= ram_a_15_0_wdata;
        ram_a_15_0_rdata_out <= ram_a_15_0_wdata;
      end else begin
        ram_a_15_0_rdata_out <= mem[ram_a_15_0_addr];
      end
    end 
  end


endmodule



module ram_a_16
(
  input CLK,
  input [20-1:0] ram_a_16_0_addr,
  output [32-1:0] ram_a_16_0_rdata,
  input [32-1:0] ram_a_16_0_wdata,
  input ram_a_16_0_wenable,
  input ram_a_16_0_enable
);

  reg [32-1:0] ram_a_16_0_rdata_out;
  assign ram_a_16_0_rdata = ram_a_16_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_a_16_0_enable) begin
      if(ram_a_16_0_wenable) begin
        mem[ram_a_16_0_addr] <= ram_a_16_0_wdata;
        ram_a_16_0_rdata_out <= ram_a_16_0_wdata;
      end else begin
        ram_a_16_0_rdata_out <= mem[ram_a_16_0_addr];
      end
    end 
  end


endmodule



module ram_a_17
(
  input CLK,
  input [20-1:0] ram_a_17_0_addr,
  output [32-1:0] ram_a_17_0_rdata,
  input [32-1:0] ram_a_17_0_wdata,
  input ram_a_17_0_wenable,
  input ram_a_17_0_enable
);

  reg [32-1:0] ram_a_17_0_rdata_out;
  assign ram_a_17_0_rdata = ram_a_17_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_a_17_0_enable) begin
      if(ram_a_17_0_wenable) begin
        mem[ram_a_17_0_addr] <= ram_a_17_0_wdata;
        ram_a_17_0_rdata_out <= ram_a_17_0_wdata;
      end else begin
        ram_a_17_0_rdata_out <= mem[ram_a_17_0_addr];
      end
    end 
  end


endmodule



module ram_a_18
(
  input CLK,
  input [20-1:0] ram_a_18_0_addr,
  output [32-1:0] ram_a_18_0_rdata,
  input [32-1:0] ram_a_18_0_wdata,
  input ram_a_18_0_wenable,
  input ram_a_18_0_enable
);

  reg [32-1:0] ram_a_18_0_rdata_out;
  assign ram_a_18_0_rdata = ram_a_18_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_a_18_0_enable) begin
      if(ram_a_18_0_wenable) begin
        mem[ram_a_18_0_addr] <= ram_a_18_0_wdata;
        ram_a_18_0_rdata_out <= ram_a_18_0_wdata;
      end else begin
        ram_a_18_0_rdata_out <= mem[ram_a_18_0_addr];
      end
    end 
  end


endmodule



module ram_a_19
(
  input CLK,
  input [20-1:0] ram_a_19_0_addr,
  output [32-1:0] ram_a_19_0_rdata,
  input [32-1:0] ram_a_19_0_wdata,
  input ram_a_19_0_wenable,
  input ram_a_19_0_enable
);

  reg [32-1:0] ram_a_19_0_rdata_out;
  assign ram_a_19_0_rdata = ram_a_19_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_a_19_0_enable) begin
      if(ram_a_19_0_wenable) begin
        mem[ram_a_19_0_addr] <= ram_a_19_0_wdata;
        ram_a_19_0_rdata_out <= ram_a_19_0_wdata;
      end else begin
        ram_a_19_0_rdata_out <= mem[ram_a_19_0_addr];
      end
    end 
  end


endmodule



module ram_a_20
(
  input CLK,
  input [20-1:0] ram_a_20_0_addr,
  output [32-1:0] ram_a_20_0_rdata,
  input [32-1:0] ram_a_20_0_wdata,
  input ram_a_20_0_wenable,
  input ram_a_20_0_enable
);

  reg [32-1:0] ram_a_20_0_rdata_out;
  assign ram_a_20_0_rdata = ram_a_20_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_a_20_0_enable) begin
      if(ram_a_20_0_wenable) begin
        mem[ram_a_20_0_addr] <= ram_a_20_0_wdata;
        ram_a_20_0_rdata_out <= ram_a_20_0_wdata;
      end else begin
        ram_a_20_0_rdata_out <= mem[ram_a_20_0_addr];
      end
    end 
  end


endmodule



module ram_a_21
(
  input CLK,
  input [20-1:0] ram_a_21_0_addr,
  output [32-1:0] ram_a_21_0_rdata,
  input [32-1:0] ram_a_21_0_wdata,
  input ram_a_21_0_wenable,
  input ram_a_21_0_enable
);

  reg [32-1:0] ram_a_21_0_rdata_out;
  assign ram_a_21_0_rdata = ram_a_21_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_a_21_0_enable) begin
      if(ram_a_21_0_wenable) begin
        mem[ram_a_21_0_addr] <= ram_a_21_0_wdata;
        ram_a_21_0_rdata_out <= ram_a_21_0_wdata;
      end else begin
        ram_a_21_0_rdata_out <= mem[ram_a_21_0_addr];
      end
    end 
  end


endmodule



module ram_a_22
(
  input CLK,
  input [20-1:0] ram_a_22_0_addr,
  output [32-1:0] ram_a_22_0_rdata,
  input [32-1:0] ram_a_22_0_wdata,
  input ram_a_22_0_wenable,
  input ram_a_22_0_enable
);

  reg [32-1:0] ram_a_22_0_rdata_out;
  assign ram_a_22_0_rdata = ram_a_22_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_a_22_0_enable) begin
      if(ram_a_22_0_wenable) begin
        mem[ram_a_22_0_addr] <= ram_a_22_0_wdata;
        ram_a_22_0_rdata_out <= ram_a_22_0_wdata;
      end else begin
        ram_a_22_0_rdata_out <= mem[ram_a_22_0_addr];
      end
    end 
  end


endmodule



module ram_a_23
(
  input CLK,
  input [20-1:0] ram_a_23_0_addr,
  output [32-1:0] ram_a_23_0_rdata,
  input [32-1:0] ram_a_23_0_wdata,
  input ram_a_23_0_wenable,
  input ram_a_23_0_enable
);

  reg [32-1:0] ram_a_23_0_rdata_out;
  assign ram_a_23_0_rdata = ram_a_23_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_a_23_0_enable) begin
      if(ram_a_23_0_wenable) begin
        mem[ram_a_23_0_addr] <= ram_a_23_0_wdata;
        ram_a_23_0_rdata_out <= ram_a_23_0_wdata;
      end else begin
        ram_a_23_0_rdata_out <= mem[ram_a_23_0_addr];
      end
    end 
  end


endmodule



module ram_a_24
(
  input CLK,
  input [20-1:0] ram_a_24_0_addr,
  output [32-1:0] ram_a_24_0_rdata,
  input [32-1:0] ram_a_24_0_wdata,
  input ram_a_24_0_wenable,
  input ram_a_24_0_enable
);

  reg [32-1:0] ram_a_24_0_rdata_out;
  assign ram_a_24_0_rdata = ram_a_24_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_a_24_0_enable) begin
      if(ram_a_24_0_wenable) begin
        mem[ram_a_24_0_addr] <= ram_a_24_0_wdata;
        ram_a_24_0_rdata_out <= ram_a_24_0_wdata;
      end else begin
        ram_a_24_0_rdata_out <= mem[ram_a_24_0_addr];
      end
    end 
  end


endmodule



module ram_a_25
(
  input CLK,
  input [20-1:0] ram_a_25_0_addr,
  output [32-1:0] ram_a_25_0_rdata,
  input [32-1:0] ram_a_25_0_wdata,
  input ram_a_25_0_wenable,
  input ram_a_25_0_enable
);

  reg [32-1:0] ram_a_25_0_rdata_out;
  assign ram_a_25_0_rdata = ram_a_25_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_a_25_0_enable) begin
      if(ram_a_25_0_wenable) begin
        mem[ram_a_25_0_addr] <= ram_a_25_0_wdata;
        ram_a_25_0_rdata_out <= ram_a_25_0_wdata;
      end else begin
        ram_a_25_0_rdata_out <= mem[ram_a_25_0_addr];
      end
    end 
  end


endmodule



module ram_a_26
(
  input CLK,
  input [20-1:0] ram_a_26_0_addr,
  output [32-1:0] ram_a_26_0_rdata,
  input [32-1:0] ram_a_26_0_wdata,
  input ram_a_26_0_wenable,
  input ram_a_26_0_enable
);

  reg [32-1:0] ram_a_26_0_rdata_out;
  assign ram_a_26_0_rdata = ram_a_26_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_a_26_0_enable) begin
      if(ram_a_26_0_wenable) begin
        mem[ram_a_26_0_addr] <= ram_a_26_0_wdata;
        ram_a_26_0_rdata_out <= ram_a_26_0_wdata;
      end else begin
        ram_a_26_0_rdata_out <= mem[ram_a_26_0_addr];
      end
    end 
  end


endmodule



module ram_a_27
(
  input CLK,
  input [20-1:0] ram_a_27_0_addr,
  output [32-1:0] ram_a_27_0_rdata,
  input [32-1:0] ram_a_27_0_wdata,
  input ram_a_27_0_wenable,
  input ram_a_27_0_enable
);

  reg [32-1:0] ram_a_27_0_rdata_out;
  assign ram_a_27_0_rdata = ram_a_27_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_a_27_0_enable) begin
      if(ram_a_27_0_wenable) begin
        mem[ram_a_27_0_addr] <= ram_a_27_0_wdata;
        ram_a_27_0_rdata_out <= ram_a_27_0_wdata;
      end else begin
        ram_a_27_0_rdata_out <= mem[ram_a_27_0_addr];
      end
    end 
  end


endmodule



module ram_a_28
(
  input CLK,
  input [20-1:0] ram_a_28_0_addr,
  output [32-1:0] ram_a_28_0_rdata,
  input [32-1:0] ram_a_28_0_wdata,
  input ram_a_28_0_wenable,
  input ram_a_28_0_enable
);

  reg [32-1:0] ram_a_28_0_rdata_out;
  assign ram_a_28_0_rdata = ram_a_28_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_a_28_0_enable) begin
      if(ram_a_28_0_wenable) begin
        mem[ram_a_28_0_addr] <= ram_a_28_0_wdata;
        ram_a_28_0_rdata_out <= ram_a_28_0_wdata;
      end else begin
        ram_a_28_0_rdata_out <= mem[ram_a_28_0_addr];
      end
    end 
  end


endmodule



module ram_a_29
(
  input CLK,
  input [20-1:0] ram_a_29_0_addr,
  output [32-1:0] ram_a_29_0_rdata,
  input [32-1:0] ram_a_29_0_wdata,
  input ram_a_29_0_wenable,
  input ram_a_29_0_enable
);

  reg [32-1:0] ram_a_29_0_rdata_out;
  assign ram_a_29_0_rdata = ram_a_29_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_a_29_0_enable) begin
      if(ram_a_29_0_wenable) begin
        mem[ram_a_29_0_addr] <= ram_a_29_0_wdata;
        ram_a_29_0_rdata_out <= ram_a_29_0_wdata;
      end else begin
        ram_a_29_0_rdata_out <= mem[ram_a_29_0_addr];
      end
    end 
  end


endmodule



module ram_a_30
(
  input CLK,
  input [20-1:0] ram_a_30_0_addr,
  output [32-1:0] ram_a_30_0_rdata,
  input [32-1:0] ram_a_30_0_wdata,
  input ram_a_30_0_wenable,
  input ram_a_30_0_enable
);

  reg [32-1:0] ram_a_30_0_rdata_out;
  assign ram_a_30_0_rdata = ram_a_30_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_a_30_0_enable) begin
      if(ram_a_30_0_wenable) begin
        mem[ram_a_30_0_addr] <= ram_a_30_0_wdata;
        ram_a_30_0_rdata_out <= ram_a_30_0_wdata;
      end else begin
        ram_a_30_0_rdata_out <= mem[ram_a_30_0_addr];
      end
    end 
  end


endmodule



module ram_a_31
(
  input CLK,
  input [20-1:0] ram_a_31_0_addr,
  output [32-1:0] ram_a_31_0_rdata,
  input [32-1:0] ram_a_31_0_wdata,
  input ram_a_31_0_wenable,
  input ram_a_31_0_enable
);

  reg [32-1:0] ram_a_31_0_rdata_out;
  assign ram_a_31_0_rdata = ram_a_31_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_a_31_0_enable) begin
      if(ram_a_31_0_wenable) begin
        mem[ram_a_31_0_addr] <= ram_a_31_0_wdata;
        ram_a_31_0_rdata_out <= ram_a_31_0_wdata;
      end else begin
        ram_a_31_0_rdata_out <= mem[ram_a_31_0_addr];
      end
    end 
  end


endmodule



module ram_b_0
(
  input CLK,
  input [20-1:0] ram_b_0_0_addr,
  output [32-1:0] ram_b_0_0_rdata,
  input [32-1:0] ram_b_0_0_wdata,
  input ram_b_0_0_wenable,
  input ram_b_0_0_enable
);

  reg [32-1:0] ram_b_0_0_rdata_out;
  assign ram_b_0_0_rdata = ram_b_0_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_b_0_0_enable) begin
      if(ram_b_0_0_wenable) begin
        mem[ram_b_0_0_addr] <= ram_b_0_0_wdata;
        ram_b_0_0_rdata_out <= ram_b_0_0_wdata;
      end else begin
        ram_b_0_0_rdata_out <= mem[ram_b_0_0_addr];
      end
    end 
  end


endmodule



module ram_b_1
(
  input CLK,
  input [20-1:0] ram_b_1_0_addr,
  output [32-1:0] ram_b_1_0_rdata,
  input [32-1:0] ram_b_1_0_wdata,
  input ram_b_1_0_wenable,
  input ram_b_1_0_enable
);

  reg [32-1:0] ram_b_1_0_rdata_out;
  assign ram_b_1_0_rdata = ram_b_1_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_b_1_0_enable) begin
      if(ram_b_1_0_wenable) begin
        mem[ram_b_1_0_addr] <= ram_b_1_0_wdata;
        ram_b_1_0_rdata_out <= ram_b_1_0_wdata;
      end else begin
        ram_b_1_0_rdata_out <= mem[ram_b_1_0_addr];
      end
    end 
  end


endmodule



module ram_b_2
(
  input CLK,
  input [20-1:0] ram_b_2_0_addr,
  output [32-1:0] ram_b_2_0_rdata,
  input [32-1:0] ram_b_2_0_wdata,
  input ram_b_2_0_wenable,
  input ram_b_2_0_enable
);

  reg [32-1:0] ram_b_2_0_rdata_out;
  assign ram_b_2_0_rdata = ram_b_2_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_b_2_0_enable) begin
      if(ram_b_2_0_wenable) begin
        mem[ram_b_2_0_addr] <= ram_b_2_0_wdata;
        ram_b_2_0_rdata_out <= ram_b_2_0_wdata;
      end else begin
        ram_b_2_0_rdata_out <= mem[ram_b_2_0_addr];
      end
    end 
  end


endmodule



module ram_b_3
(
  input CLK,
  input [20-1:0] ram_b_3_0_addr,
  output [32-1:0] ram_b_3_0_rdata,
  input [32-1:0] ram_b_3_0_wdata,
  input ram_b_3_0_wenable,
  input ram_b_3_0_enable
);

  reg [32-1:0] ram_b_3_0_rdata_out;
  assign ram_b_3_0_rdata = ram_b_3_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_b_3_0_enable) begin
      if(ram_b_3_0_wenable) begin
        mem[ram_b_3_0_addr] <= ram_b_3_0_wdata;
        ram_b_3_0_rdata_out <= ram_b_3_0_wdata;
      end else begin
        ram_b_3_0_rdata_out <= mem[ram_b_3_0_addr];
      end
    end 
  end


endmodule



module ram_b_4
(
  input CLK,
  input [20-1:0] ram_b_4_0_addr,
  output [32-1:0] ram_b_4_0_rdata,
  input [32-1:0] ram_b_4_0_wdata,
  input ram_b_4_0_wenable,
  input ram_b_4_0_enable
);

  reg [32-1:0] ram_b_4_0_rdata_out;
  assign ram_b_4_0_rdata = ram_b_4_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_b_4_0_enable) begin
      if(ram_b_4_0_wenable) begin
        mem[ram_b_4_0_addr] <= ram_b_4_0_wdata;
        ram_b_4_0_rdata_out <= ram_b_4_0_wdata;
      end else begin
        ram_b_4_0_rdata_out <= mem[ram_b_4_0_addr];
      end
    end 
  end


endmodule



module ram_b_5
(
  input CLK,
  input [20-1:0] ram_b_5_0_addr,
  output [32-1:0] ram_b_5_0_rdata,
  input [32-1:0] ram_b_5_0_wdata,
  input ram_b_5_0_wenable,
  input ram_b_5_0_enable
);

  reg [32-1:0] ram_b_5_0_rdata_out;
  assign ram_b_5_0_rdata = ram_b_5_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_b_5_0_enable) begin
      if(ram_b_5_0_wenable) begin
        mem[ram_b_5_0_addr] <= ram_b_5_0_wdata;
        ram_b_5_0_rdata_out <= ram_b_5_0_wdata;
      end else begin
        ram_b_5_0_rdata_out <= mem[ram_b_5_0_addr];
      end
    end 
  end


endmodule



module ram_b_6
(
  input CLK,
  input [20-1:0] ram_b_6_0_addr,
  output [32-1:0] ram_b_6_0_rdata,
  input [32-1:0] ram_b_6_0_wdata,
  input ram_b_6_0_wenable,
  input ram_b_6_0_enable
);

  reg [32-1:0] ram_b_6_0_rdata_out;
  assign ram_b_6_0_rdata = ram_b_6_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_b_6_0_enable) begin
      if(ram_b_6_0_wenable) begin
        mem[ram_b_6_0_addr] <= ram_b_6_0_wdata;
        ram_b_6_0_rdata_out <= ram_b_6_0_wdata;
      end else begin
        ram_b_6_0_rdata_out <= mem[ram_b_6_0_addr];
      end
    end 
  end


endmodule



module ram_b_7
(
  input CLK,
  input [20-1:0] ram_b_7_0_addr,
  output [32-1:0] ram_b_7_0_rdata,
  input [32-1:0] ram_b_7_0_wdata,
  input ram_b_7_0_wenable,
  input ram_b_7_0_enable
);

  reg [32-1:0] ram_b_7_0_rdata_out;
  assign ram_b_7_0_rdata = ram_b_7_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_b_7_0_enable) begin
      if(ram_b_7_0_wenable) begin
        mem[ram_b_7_0_addr] <= ram_b_7_0_wdata;
        ram_b_7_0_rdata_out <= ram_b_7_0_wdata;
      end else begin
        ram_b_7_0_rdata_out <= mem[ram_b_7_0_addr];
      end
    end 
  end


endmodule



module ram_b_8
(
  input CLK,
  input [20-1:0] ram_b_8_0_addr,
  output [32-1:0] ram_b_8_0_rdata,
  input [32-1:0] ram_b_8_0_wdata,
  input ram_b_8_0_wenable,
  input ram_b_8_0_enable
);

  reg [32-1:0] ram_b_8_0_rdata_out;
  assign ram_b_8_0_rdata = ram_b_8_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_b_8_0_enable) begin
      if(ram_b_8_0_wenable) begin
        mem[ram_b_8_0_addr] <= ram_b_8_0_wdata;
        ram_b_8_0_rdata_out <= ram_b_8_0_wdata;
      end else begin
        ram_b_8_0_rdata_out <= mem[ram_b_8_0_addr];
      end
    end 
  end


endmodule



module ram_b_9
(
  input CLK,
  input [20-1:0] ram_b_9_0_addr,
  output [32-1:0] ram_b_9_0_rdata,
  input [32-1:0] ram_b_9_0_wdata,
  input ram_b_9_0_wenable,
  input ram_b_9_0_enable
);

  reg [32-1:0] ram_b_9_0_rdata_out;
  assign ram_b_9_0_rdata = ram_b_9_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_b_9_0_enable) begin
      if(ram_b_9_0_wenable) begin
        mem[ram_b_9_0_addr] <= ram_b_9_0_wdata;
        ram_b_9_0_rdata_out <= ram_b_9_0_wdata;
      end else begin
        ram_b_9_0_rdata_out <= mem[ram_b_9_0_addr];
      end
    end 
  end


endmodule



module ram_b_10
(
  input CLK,
  input [20-1:0] ram_b_10_0_addr,
  output [32-1:0] ram_b_10_0_rdata,
  input [32-1:0] ram_b_10_0_wdata,
  input ram_b_10_0_wenable,
  input ram_b_10_0_enable
);

  reg [32-1:0] ram_b_10_0_rdata_out;
  assign ram_b_10_0_rdata = ram_b_10_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_b_10_0_enable) begin
      if(ram_b_10_0_wenable) begin
        mem[ram_b_10_0_addr] <= ram_b_10_0_wdata;
        ram_b_10_0_rdata_out <= ram_b_10_0_wdata;
      end else begin
        ram_b_10_0_rdata_out <= mem[ram_b_10_0_addr];
      end
    end 
  end


endmodule



module ram_b_11
(
  input CLK,
  input [20-1:0] ram_b_11_0_addr,
  output [32-1:0] ram_b_11_0_rdata,
  input [32-1:0] ram_b_11_0_wdata,
  input ram_b_11_0_wenable,
  input ram_b_11_0_enable
);

  reg [32-1:0] ram_b_11_0_rdata_out;
  assign ram_b_11_0_rdata = ram_b_11_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_b_11_0_enable) begin
      if(ram_b_11_0_wenable) begin
        mem[ram_b_11_0_addr] <= ram_b_11_0_wdata;
        ram_b_11_0_rdata_out <= ram_b_11_0_wdata;
      end else begin
        ram_b_11_0_rdata_out <= mem[ram_b_11_0_addr];
      end
    end 
  end


endmodule



module ram_b_12
(
  input CLK,
  input [20-1:0] ram_b_12_0_addr,
  output [32-1:0] ram_b_12_0_rdata,
  input [32-1:0] ram_b_12_0_wdata,
  input ram_b_12_0_wenable,
  input ram_b_12_0_enable
);

  reg [32-1:0] ram_b_12_0_rdata_out;
  assign ram_b_12_0_rdata = ram_b_12_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_b_12_0_enable) begin
      if(ram_b_12_0_wenable) begin
        mem[ram_b_12_0_addr] <= ram_b_12_0_wdata;
        ram_b_12_0_rdata_out <= ram_b_12_0_wdata;
      end else begin
        ram_b_12_0_rdata_out <= mem[ram_b_12_0_addr];
      end
    end 
  end


endmodule



module ram_b_13
(
  input CLK,
  input [20-1:0] ram_b_13_0_addr,
  output [32-1:0] ram_b_13_0_rdata,
  input [32-1:0] ram_b_13_0_wdata,
  input ram_b_13_0_wenable,
  input ram_b_13_0_enable
);

  reg [32-1:0] ram_b_13_0_rdata_out;
  assign ram_b_13_0_rdata = ram_b_13_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_b_13_0_enable) begin
      if(ram_b_13_0_wenable) begin
        mem[ram_b_13_0_addr] <= ram_b_13_0_wdata;
        ram_b_13_0_rdata_out <= ram_b_13_0_wdata;
      end else begin
        ram_b_13_0_rdata_out <= mem[ram_b_13_0_addr];
      end
    end 
  end


endmodule



module ram_b_14
(
  input CLK,
  input [20-1:0] ram_b_14_0_addr,
  output [32-1:0] ram_b_14_0_rdata,
  input [32-1:0] ram_b_14_0_wdata,
  input ram_b_14_0_wenable,
  input ram_b_14_0_enable
);

  reg [32-1:0] ram_b_14_0_rdata_out;
  assign ram_b_14_0_rdata = ram_b_14_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_b_14_0_enable) begin
      if(ram_b_14_0_wenable) begin
        mem[ram_b_14_0_addr] <= ram_b_14_0_wdata;
        ram_b_14_0_rdata_out <= ram_b_14_0_wdata;
      end else begin
        ram_b_14_0_rdata_out <= mem[ram_b_14_0_addr];
      end
    end 
  end


endmodule



module ram_b_15
(
  input CLK,
  input [20-1:0] ram_b_15_0_addr,
  output [32-1:0] ram_b_15_0_rdata,
  input [32-1:0] ram_b_15_0_wdata,
  input ram_b_15_0_wenable,
  input ram_b_15_0_enable
);

  reg [32-1:0] ram_b_15_0_rdata_out;
  assign ram_b_15_0_rdata = ram_b_15_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_b_15_0_enable) begin
      if(ram_b_15_0_wenable) begin
        mem[ram_b_15_0_addr] <= ram_b_15_0_wdata;
        ram_b_15_0_rdata_out <= ram_b_15_0_wdata;
      end else begin
        ram_b_15_0_rdata_out <= mem[ram_b_15_0_addr];
      end
    end 
  end


endmodule



module ram_b_16
(
  input CLK,
  input [20-1:0] ram_b_16_0_addr,
  output [32-1:0] ram_b_16_0_rdata,
  input [32-1:0] ram_b_16_0_wdata,
  input ram_b_16_0_wenable,
  input ram_b_16_0_enable
);

  reg [32-1:0] ram_b_16_0_rdata_out;
  assign ram_b_16_0_rdata = ram_b_16_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_b_16_0_enable) begin
      if(ram_b_16_0_wenable) begin
        mem[ram_b_16_0_addr] <= ram_b_16_0_wdata;
        ram_b_16_0_rdata_out <= ram_b_16_0_wdata;
      end else begin
        ram_b_16_0_rdata_out <= mem[ram_b_16_0_addr];
      end
    end 
  end


endmodule



module ram_b_17
(
  input CLK,
  input [20-1:0] ram_b_17_0_addr,
  output [32-1:0] ram_b_17_0_rdata,
  input [32-1:0] ram_b_17_0_wdata,
  input ram_b_17_0_wenable,
  input ram_b_17_0_enable
);

  reg [32-1:0] ram_b_17_0_rdata_out;
  assign ram_b_17_0_rdata = ram_b_17_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_b_17_0_enable) begin
      if(ram_b_17_0_wenable) begin
        mem[ram_b_17_0_addr] <= ram_b_17_0_wdata;
        ram_b_17_0_rdata_out <= ram_b_17_0_wdata;
      end else begin
        ram_b_17_0_rdata_out <= mem[ram_b_17_0_addr];
      end
    end 
  end


endmodule



module ram_b_18
(
  input CLK,
  input [20-1:0] ram_b_18_0_addr,
  output [32-1:0] ram_b_18_0_rdata,
  input [32-1:0] ram_b_18_0_wdata,
  input ram_b_18_0_wenable,
  input ram_b_18_0_enable
);

  reg [32-1:0] ram_b_18_0_rdata_out;
  assign ram_b_18_0_rdata = ram_b_18_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_b_18_0_enable) begin
      if(ram_b_18_0_wenable) begin
        mem[ram_b_18_0_addr] <= ram_b_18_0_wdata;
        ram_b_18_0_rdata_out <= ram_b_18_0_wdata;
      end else begin
        ram_b_18_0_rdata_out <= mem[ram_b_18_0_addr];
      end
    end 
  end


endmodule



module ram_b_19
(
  input CLK,
  input [20-1:0] ram_b_19_0_addr,
  output [32-1:0] ram_b_19_0_rdata,
  input [32-1:0] ram_b_19_0_wdata,
  input ram_b_19_0_wenable,
  input ram_b_19_0_enable
);

  reg [32-1:0] ram_b_19_0_rdata_out;
  assign ram_b_19_0_rdata = ram_b_19_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_b_19_0_enable) begin
      if(ram_b_19_0_wenable) begin
        mem[ram_b_19_0_addr] <= ram_b_19_0_wdata;
        ram_b_19_0_rdata_out <= ram_b_19_0_wdata;
      end else begin
        ram_b_19_0_rdata_out <= mem[ram_b_19_0_addr];
      end
    end 
  end


endmodule



module ram_b_20
(
  input CLK,
  input [20-1:0] ram_b_20_0_addr,
  output [32-1:0] ram_b_20_0_rdata,
  input [32-1:0] ram_b_20_0_wdata,
  input ram_b_20_0_wenable,
  input ram_b_20_0_enable
);

  reg [32-1:0] ram_b_20_0_rdata_out;
  assign ram_b_20_0_rdata = ram_b_20_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_b_20_0_enable) begin
      if(ram_b_20_0_wenable) begin
        mem[ram_b_20_0_addr] <= ram_b_20_0_wdata;
        ram_b_20_0_rdata_out <= ram_b_20_0_wdata;
      end else begin
        ram_b_20_0_rdata_out <= mem[ram_b_20_0_addr];
      end
    end 
  end


endmodule



module ram_b_21
(
  input CLK,
  input [20-1:0] ram_b_21_0_addr,
  output [32-1:0] ram_b_21_0_rdata,
  input [32-1:0] ram_b_21_0_wdata,
  input ram_b_21_0_wenable,
  input ram_b_21_0_enable
);

  reg [32-1:0] ram_b_21_0_rdata_out;
  assign ram_b_21_0_rdata = ram_b_21_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_b_21_0_enable) begin
      if(ram_b_21_0_wenable) begin
        mem[ram_b_21_0_addr] <= ram_b_21_0_wdata;
        ram_b_21_0_rdata_out <= ram_b_21_0_wdata;
      end else begin
        ram_b_21_0_rdata_out <= mem[ram_b_21_0_addr];
      end
    end 
  end


endmodule



module ram_b_22
(
  input CLK,
  input [20-1:0] ram_b_22_0_addr,
  output [32-1:0] ram_b_22_0_rdata,
  input [32-1:0] ram_b_22_0_wdata,
  input ram_b_22_0_wenable,
  input ram_b_22_0_enable
);

  reg [32-1:0] ram_b_22_0_rdata_out;
  assign ram_b_22_0_rdata = ram_b_22_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_b_22_0_enable) begin
      if(ram_b_22_0_wenable) begin
        mem[ram_b_22_0_addr] <= ram_b_22_0_wdata;
        ram_b_22_0_rdata_out <= ram_b_22_0_wdata;
      end else begin
        ram_b_22_0_rdata_out <= mem[ram_b_22_0_addr];
      end
    end 
  end


endmodule



module ram_b_23
(
  input CLK,
  input [20-1:0] ram_b_23_0_addr,
  output [32-1:0] ram_b_23_0_rdata,
  input [32-1:0] ram_b_23_0_wdata,
  input ram_b_23_0_wenable,
  input ram_b_23_0_enable
);

  reg [32-1:0] ram_b_23_0_rdata_out;
  assign ram_b_23_0_rdata = ram_b_23_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_b_23_0_enable) begin
      if(ram_b_23_0_wenable) begin
        mem[ram_b_23_0_addr] <= ram_b_23_0_wdata;
        ram_b_23_0_rdata_out <= ram_b_23_0_wdata;
      end else begin
        ram_b_23_0_rdata_out <= mem[ram_b_23_0_addr];
      end
    end 
  end


endmodule



module ram_b_24
(
  input CLK,
  input [20-1:0] ram_b_24_0_addr,
  output [32-1:0] ram_b_24_0_rdata,
  input [32-1:0] ram_b_24_0_wdata,
  input ram_b_24_0_wenable,
  input ram_b_24_0_enable
);

  reg [32-1:0] ram_b_24_0_rdata_out;
  assign ram_b_24_0_rdata = ram_b_24_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_b_24_0_enable) begin
      if(ram_b_24_0_wenable) begin
        mem[ram_b_24_0_addr] <= ram_b_24_0_wdata;
        ram_b_24_0_rdata_out <= ram_b_24_0_wdata;
      end else begin
        ram_b_24_0_rdata_out <= mem[ram_b_24_0_addr];
      end
    end 
  end


endmodule



module ram_b_25
(
  input CLK,
  input [20-1:0] ram_b_25_0_addr,
  output [32-1:0] ram_b_25_0_rdata,
  input [32-1:0] ram_b_25_0_wdata,
  input ram_b_25_0_wenable,
  input ram_b_25_0_enable
);

  reg [32-1:0] ram_b_25_0_rdata_out;
  assign ram_b_25_0_rdata = ram_b_25_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_b_25_0_enable) begin
      if(ram_b_25_0_wenable) begin
        mem[ram_b_25_0_addr] <= ram_b_25_0_wdata;
        ram_b_25_0_rdata_out <= ram_b_25_0_wdata;
      end else begin
        ram_b_25_0_rdata_out <= mem[ram_b_25_0_addr];
      end
    end 
  end


endmodule



module ram_b_26
(
  input CLK,
  input [20-1:0] ram_b_26_0_addr,
  output [32-1:0] ram_b_26_0_rdata,
  input [32-1:0] ram_b_26_0_wdata,
  input ram_b_26_0_wenable,
  input ram_b_26_0_enable
);

  reg [32-1:0] ram_b_26_0_rdata_out;
  assign ram_b_26_0_rdata = ram_b_26_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_b_26_0_enable) begin
      if(ram_b_26_0_wenable) begin
        mem[ram_b_26_0_addr] <= ram_b_26_0_wdata;
        ram_b_26_0_rdata_out <= ram_b_26_0_wdata;
      end else begin
        ram_b_26_0_rdata_out <= mem[ram_b_26_0_addr];
      end
    end 
  end


endmodule



module ram_b_27
(
  input CLK,
  input [20-1:0] ram_b_27_0_addr,
  output [32-1:0] ram_b_27_0_rdata,
  input [32-1:0] ram_b_27_0_wdata,
  input ram_b_27_0_wenable,
  input ram_b_27_0_enable
);

  reg [32-1:0] ram_b_27_0_rdata_out;
  assign ram_b_27_0_rdata = ram_b_27_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_b_27_0_enable) begin
      if(ram_b_27_0_wenable) begin
        mem[ram_b_27_0_addr] <= ram_b_27_0_wdata;
        ram_b_27_0_rdata_out <= ram_b_27_0_wdata;
      end else begin
        ram_b_27_0_rdata_out <= mem[ram_b_27_0_addr];
      end
    end 
  end


endmodule



module ram_b_28
(
  input CLK,
  input [20-1:0] ram_b_28_0_addr,
  output [32-1:0] ram_b_28_0_rdata,
  input [32-1:0] ram_b_28_0_wdata,
  input ram_b_28_0_wenable,
  input ram_b_28_0_enable
);

  reg [32-1:0] ram_b_28_0_rdata_out;
  assign ram_b_28_0_rdata = ram_b_28_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_b_28_0_enable) begin
      if(ram_b_28_0_wenable) begin
        mem[ram_b_28_0_addr] <= ram_b_28_0_wdata;
        ram_b_28_0_rdata_out <= ram_b_28_0_wdata;
      end else begin
        ram_b_28_0_rdata_out <= mem[ram_b_28_0_addr];
      end
    end 
  end


endmodule



module ram_b_29
(
  input CLK,
  input [20-1:0] ram_b_29_0_addr,
  output [32-1:0] ram_b_29_0_rdata,
  input [32-1:0] ram_b_29_0_wdata,
  input ram_b_29_0_wenable,
  input ram_b_29_0_enable
);

  reg [32-1:0] ram_b_29_0_rdata_out;
  assign ram_b_29_0_rdata = ram_b_29_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_b_29_0_enable) begin
      if(ram_b_29_0_wenable) begin
        mem[ram_b_29_0_addr] <= ram_b_29_0_wdata;
        ram_b_29_0_rdata_out <= ram_b_29_0_wdata;
      end else begin
        ram_b_29_0_rdata_out <= mem[ram_b_29_0_addr];
      end
    end 
  end


endmodule



module ram_b_30
(
  input CLK,
  input [20-1:0] ram_b_30_0_addr,
  output [32-1:0] ram_b_30_0_rdata,
  input [32-1:0] ram_b_30_0_wdata,
  input ram_b_30_0_wenable,
  input ram_b_30_0_enable
);

  reg [32-1:0] ram_b_30_0_rdata_out;
  assign ram_b_30_0_rdata = ram_b_30_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_b_30_0_enable) begin
      if(ram_b_30_0_wenable) begin
        mem[ram_b_30_0_addr] <= ram_b_30_0_wdata;
        ram_b_30_0_rdata_out <= ram_b_30_0_wdata;
      end else begin
        ram_b_30_0_rdata_out <= mem[ram_b_30_0_addr];
      end
    end 
  end


endmodule



module ram_b_31
(
  input CLK,
  input [20-1:0] ram_b_31_0_addr,
  output [32-1:0] ram_b_31_0_rdata,
  input [32-1:0] ram_b_31_0_wdata,
  input ram_b_31_0_wenable,
  input ram_b_31_0_enable
);

  reg [32-1:0] ram_b_31_0_rdata_out;
  assign ram_b_31_0_rdata = ram_b_31_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_b_31_0_enable) begin
      if(ram_b_31_0_wenable) begin
        mem[ram_b_31_0_addr] <= ram_b_31_0_wdata;
        ram_b_31_0_rdata_out <= ram_b_31_0_wdata;
      end else begin
        ram_b_31_0_rdata_out <= mem[ram_b_31_0_addr];
      end
    end 
  end


endmodule



module ram_c_0
(
  input CLK,
  input [20-1:0] ram_c_0_0_addr,
  output [32-1:0] ram_c_0_0_rdata,
  input [32-1:0] ram_c_0_0_wdata,
  input ram_c_0_0_wenable,
  input ram_c_0_0_enable
);

  reg [32-1:0] ram_c_0_0_rdata_out;
  assign ram_c_0_0_rdata = ram_c_0_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_c_0_0_enable) begin
      if(ram_c_0_0_wenable) begin
        mem[ram_c_0_0_addr] <= ram_c_0_0_wdata;
        ram_c_0_0_rdata_out <= ram_c_0_0_wdata;
      end else begin
        ram_c_0_0_rdata_out <= mem[ram_c_0_0_addr];
      end
    end 
  end


endmodule



module ram_c_1
(
  input CLK,
  input [20-1:0] ram_c_1_0_addr,
  output [32-1:0] ram_c_1_0_rdata,
  input [32-1:0] ram_c_1_0_wdata,
  input ram_c_1_0_wenable,
  input ram_c_1_0_enable
);

  reg [32-1:0] ram_c_1_0_rdata_out;
  assign ram_c_1_0_rdata = ram_c_1_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_c_1_0_enable) begin
      if(ram_c_1_0_wenable) begin
        mem[ram_c_1_0_addr] <= ram_c_1_0_wdata;
        ram_c_1_0_rdata_out <= ram_c_1_0_wdata;
      end else begin
        ram_c_1_0_rdata_out <= mem[ram_c_1_0_addr];
      end
    end 
  end


endmodule



module ram_c_2
(
  input CLK,
  input [20-1:0] ram_c_2_0_addr,
  output [32-1:0] ram_c_2_0_rdata,
  input [32-1:0] ram_c_2_0_wdata,
  input ram_c_2_0_wenable,
  input ram_c_2_0_enable
);

  reg [32-1:0] ram_c_2_0_rdata_out;
  assign ram_c_2_0_rdata = ram_c_2_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_c_2_0_enable) begin
      if(ram_c_2_0_wenable) begin
        mem[ram_c_2_0_addr] <= ram_c_2_0_wdata;
        ram_c_2_0_rdata_out <= ram_c_2_0_wdata;
      end else begin
        ram_c_2_0_rdata_out <= mem[ram_c_2_0_addr];
      end
    end 
  end


endmodule



module ram_c_3
(
  input CLK,
  input [20-1:0] ram_c_3_0_addr,
  output [32-1:0] ram_c_3_0_rdata,
  input [32-1:0] ram_c_3_0_wdata,
  input ram_c_3_0_wenable,
  input ram_c_3_0_enable
);

  reg [32-1:0] ram_c_3_0_rdata_out;
  assign ram_c_3_0_rdata = ram_c_3_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_c_3_0_enable) begin
      if(ram_c_3_0_wenable) begin
        mem[ram_c_3_0_addr] <= ram_c_3_0_wdata;
        ram_c_3_0_rdata_out <= ram_c_3_0_wdata;
      end else begin
        ram_c_3_0_rdata_out <= mem[ram_c_3_0_addr];
      end
    end 
  end


endmodule



module ram_c_4
(
  input CLK,
  input [20-1:0] ram_c_4_0_addr,
  output [32-1:0] ram_c_4_0_rdata,
  input [32-1:0] ram_c_4_0_wdata,
  input ram_c_4_0_wenable,
  input ram_c_4_0_enable
);

  reg [32-1:0] ram_c_4_0_rdata_out;
  assign ram_c_4_0_rdata = ram_c_4_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_c_4_0_enable) begin
      if(ram_c_4_0_wenable) begin
        mem[ram_c_4_0_addr] <= ram_c_4_0_wdata;
        ram_c_4_0_rdata_out <= ram_c_4_0_wdata;
      end else begin
        ram_c_4_0_rdata_out <= mem[ram_c_4_0_addr];
      end
    end 
  end


endmodule



module ram_c_5
(
  input CLK,
  input [20-1:0] ram_c_5_0_addr,
  output [32-1:0] ram_c_5_0_rdata,
  input [32-1:0] ram_c_5_0_wdata,
  input ram_c_5_0_wenable,
  input ram_c_5_0_enable
);

  reg [32-1:0] ram_c_5_0_rdata_out;
  assign ram_c_5_0_rdata = ram_c_5_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_c_5_0_enable) begin
      if(ram_c_5_0_wenable) begin
        mem[ram_c_5_0_addr] <= ram_c_5_0_wdata;
        ram_c_5_0_rdata_out <= ram_c_5_0_wdata;
      end else begin
        ram_c_5_0_rdata_out <= mem[ram_c_5_0_addr];
      end
    end 
  end


endmodule



module ram_c_6
(
  input CLK,
  input [20-1:0] ram_c_6_0_addr,
  output [32-1:0] ram_c_6_0_rdata,
  input [32-1:0] ram_c_6_0_wdata,
  input ram_c_6_0_wenable,
  input ram_c_6_0_enable
);

  reg [32-1:0] ram_c_6_0_rdata_out;
  assign ram_c_6_0_rdata = ram_c_6_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_c_6_0_enable) begin
      if(ram_c_6_0_wenable) begin
        mem[ram_c_6_0_addr] <= ram_c_6_0_wdata;
        ram_c_6_0_rdata_out <= ram_c_6_0_wdata;
      end else begin
        ram_c_6_0_rdata_out <= mem[ram_c_6_0_addr];
      end
    end 
  end


endmodule



module ram_c_7
(
  input CLK,
  input [20-1:0] ram_c_7_0_addr,
  output [32-1:0] ram_c_7_0_rdata,
  input [32-1:0] ram_c_7_0_wdata,
  input ram_c_7_0_wenable,
  input ram_c_7_0_enable
);

  reg [32-1:0] ram_c_7_0_rdata_out;
  assign ram_c_7_0_rdata = ram_c_7_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_c_7_0_enable) begin
      if(ram_c_7_0_wenable) begin
        mem[ram_c_7_0_addr] <= ram_c_7_0_wdata;
        ram_c_7_0_rdata_out <= ram_c_7_0_wdata;
      end else begin
        ram_c_7_0_rdata_out <= mem[ram_c_7_0_addr];
      end
    end 
  end


endmodule



module ram_c_8
(
  input CLK,
  input [20-1:0] ram_c_8_0_addr,
  output [32-1:0] ram_c_8_0_rdata,
  input [32-1:0] ram_c_8_0_wdata,
  input ram_c_8_0_wenable,
  input ram_c_8_0_enable
);

  reg [32-1:0] ram_c_8_0_rdata_out;
  assign ram_c_8_0_rdata = ram_c_8_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_c_8_0_enable) begin
      if(ram_c_8_0_wenable) begin
        mem[ram_c_8_0_addr] <= ram_c_8_0_wdata;
        ram_c_8_0_rdata_out <= ram_c_8_0_wdata;
      end else begin
        ram_c_8_0_rdata_out <= mem[ram_c_8_0_addr];
      end
    end 
  end


endmodule



module ram_c_9
(
  input CLK,
  input [20-1:0] ram_c_9_0_addr,
  output [32-1:0] ram_c_9_0_rdata,
  input [32-1:0] ram_c_9_0_wdata,
  input ram_c_9_0_wenable,
  input ram_c_9_0_enable
);

  reg [32-1:0] ram_c_9_0_rdata_out;
  assign ram_c_9_0_rdata = ram_c_9_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_c_9_0_enable) begin
      if(ram_c_9_0_wenable) begin
        mem[ram_c_9_0_addr] <= ram_c_9_0_wdata;
        ram_c_9_0_rdata_out <= ram_c_9_0_wdata;
      end else begin
        ram_c_9_0_rdata_out <= mem[ram_c_9_0_addr];
      end
    end 
  end


endmodule



module ram_c_10
(
  input CLK,
  input [20-1:0] ram_c_10_0_addr,
  output [32-1:0] ram_c_10_0_rdata,
  input [32-1:0] ram_c_10_0_wdata,
  input ram_c_10_0_wenable,
  input ram_c_10_0_enable
);

  reg [32-1:0] ram_c_10_0_rdata_out;
  assign ram_c_10_0_rdata = ram_c_10_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_c_10_0_enable) begin
      if(ram_c_10_0_wenable) begin
        mem[ram_c_10_0_addr] <= ram_c_10_0_wdata;
        ram_c_10_0_rdata_out <= ram_c_10_0_wdata;
      end else begin
        ram_c_10_0_rdata_out <= mem[ram_c_10_0_addr];
      end
    end 
  end


endmodule



module ram_c_11
(
  input CLK,
  input [20-1:0] ram_c_11_0_addr,
  output [32-1:0] ram_c_11_0_rdata,
  input [32-1:0] ram_c_11_0_wdata,
  input ram_c_11_0_wenable,
  input ram_c_11_0_enable
);

  reg [32-1:0] ram_c_11_0_rdata_out;
  assign ram_c_11_0_rdata = ram_c_11_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_c_11_0_enable) begin
      if(ram_c_11_0_wenable) begin
        mem[ram_c_11_0_addr] <= ram_c_11_0_wdata;
        ram_c_11_0_rdata_out <= ram_c_11_0_wdata;
      end else begin
        ram_c_11_0_rdata_out <= mem[ram_c_11_0_addr];
      end
    end 
  end


endmodule



module ram_c_12
(
  input CLK,
  input [20-1:0] ram_c_12_0_addr,
  output [32-1:0] ram_c_12_0_rdata,
  input [32-1:0] ram_c_12_0_wdata,
  input ram_c_12_0_wenable,
  input ram_c_12_0_enable
);

  reg [32-1:0] ram_c_12_0_rdata_out;
  assign ram_c_12_0_rdata = ram_c_12_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_c_12_0_enable) begin
      if(ram_c_12_0_wenable) begin
        mem[ram_c_12_0_addr] <= ram_c_12_0_wdata;
        ram_c_12_0_rdata_out <= ram_c_12_0_wdata;
      end else begin
        ram_c_12_0_rdata_out <= mem[ram_c_12_0_addr];
      end
    end 
  end


endmodule



module ram_c_13
(
  input CLK,
  input [20-1:0] ram_c_13_0_addr,
  output [32-1:0] ram_c_13_0_rdata,
  input [32-1:0] ram_c_13_0_wdata,
  input ram_c_13_0_wenable,
  input ram_c_13_0_enable
);

  reg [32-1:0] ram_c_13_0_rdata_out;
  assign ram_c_13_0_rdata = ram_c_13_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_c_13_0_enable) begin
      if(ram_c_13_0_wenable) begin
        mem[ram_c_13_0_addr] <= ram_c_13_0_wdata;
        ram_c_13_0_rdata_out <= ram_c_13_0_wdata;
      end else begin
        ram_c_13_0_rdata_out <= mem[ram_c_13_0_addr];
      end
    end 
  end


endmodule



module ram_c_14
(
  input CLK,
  input [20-1:0] ram_c_14_0_addr,
  output [32-1:0] ram_c_14_0_rdata,
  input [32-1:0] ram_c_14_0_wdata,
  input ram_c_14_0_wenable,
  input ram_c_14_0_enable
);

  reg [32-1:0] ram_c_14_0_rdata_out;
  assign ram_c_14_0_rdata = ram_c_14_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_c_14_0_enable) begin
      if(ram_c_14_0_wenable) begin
        mem[ram_c_14_0_addr] <= ram_c_14_0_wdata;
        ram_c_14_0_rdata_out <= ram_c_14_0_wdata;
      end else begin
        ram_c_14_0_rdata_out <= mem[ram_c_14_0_addr];
      end
    end 
  end


endmodule



module ram_c_15
(
  input CLK,
  input [20-1:0] ram_c_15_0_addr,
  output [32-1:0] ram_c_15_0_rdata,
  input [32-1:0] ram_c_15_0_wdata,
  input ram_c_15_0_wenable,
  input ram_c_15_0_enable
);

  reg [32-1:0] ram_c_15_0_rdata_out;
  assign ram_c_15_0_rdata = ram_c_15_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_c_15_0_enable) begin
      if(ram_c_15_0_wenable) begin
        mem[ram_c_15_0_addr] <= ram_c_15_0_wdata;
        ram_c_15_0_rdata_out <= ram_c_15_0_wdata;
      end else begin
        ram_c_15_0_rdata_out <= mem[ram_c_15_0_addr];
      end
    end 
  end


endmodule



module ram_c_16
(
  input CLK,
  input [20-1:0] ram_c_16_0_addr,
  output [32-1:0] ram_c_16_0_rdata,
  input [32-1:0] ram_c_16_0_wdata,
  input ram_c_16_0_wenable,
  input ram_c_16_0_enable
);

  reg [32-1:0] ram_c_16_0_rdata_out;
  assign ram_c_16_0_rdata = ram_c_16_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_c_16_0_enable) begin
      if(ram_c_16_0_wenable) begin
        mem[ram_c_16_0_addr] <= ram_c_16_0_wdata;
        ram_c_16_0_rdata_out <= ram_c_16_0_wdata;
      end else begin
        ram_c_16_0_rdata_out <= mem[ram_c_16_0_addr];
      end
    end 
  end


endmodule



module ram_c_17
(
  input CLK,
  input [20-1:0] ram_c_17_0_addr,
  output [32-1:0] ram_c_17_0_rdata,
  input [32-1:0] ram_c_17_0_wdata,
  input ram_c_17_0_wenable,
  input ram_c_17_0_enable
);

  reg [32-1:0] ram_c_17_0_rdata_out;
  assign ram_c_17_0_rdata = ram_c_17_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_c_17_0_enable) begin
      if(ram_c_17_0_wenable) begin
        mem[ram_c_17_0_addr] <= ram_c_17_0_wdata;
        ram_c_17_0_rdata_out <= ram_c_17_0_wdata;
      end else begin
        ram_c_17_0_rdata_out <= mem[ram_c_17_0_addr];
      end
    end 
  end


endmodule



module ram_c_18
(
  input CLK,
  input [20-1:0] ram_c_18_0_addr,
  output [32-1:0] ram_c_18_0_rdata,
  input [32-1:0] ram_c_18_0_wdata,
  input ram_c_18_0_wenable,
  input ram_c_18_0_enable
);

  reg [32-1:0] ram_c_18_0_rdata_out;
  assign ram_c_18_0_rdata = ram_c_18_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_c_18_0_enable) begin
      if(ram_c_18_0_wenable) begin
        mem[ram_c_18_0_addr] <= ram_c_18_0_wdata;
        ram_c_18_0_rdata_out <= ram_c_18_0_wdata;
      end else begin
        ram_c_18_0_rdata_out <= mem[ram_c_18_0_addr];
      end
    end 
  end


endmodule



module ram_c_19
(
  input CLK,
  input [20-1:0] ram_c_19_0_addr,
  output [32-1:0] ram_c_19_0_rdata,
  input [32-1:0] ram_c_19_0_wdata,
  input ram_c_19_0_wenable,
  input ram_c_19_0_enable
);

  reg [32-1:0] ram_c_19_0_rdata_out;
  assign ram_c_19_0_rdata = ram_c_19_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_c_19_0_enable) begin
      if(ram_c_19_0_wenable) begin
        mem[ram_c_19_0_addr] <= ram_c_19_0_wdata;
        ram_c_19_0_rdata_out <= ram_c_19_0_wdata;
      end else begin
        ram_c_19_0_rdata_out <= mem[ram_c_19_0_addr];
      end
    end 
  end


endmodule



module ram_c_20
(
  input CLK,
  input [20-1:0] ram_c_20_0_addr,
  output [32-1:0] ram_c_20_0_rdata,
  input [32-1:0] ram_c_20_0_wdata,
  input ram_c_20_0_wenable,
  input ram_c_20_0_enable
);

  reg [32-1:0] ram_c_20_0_rdata_out;
  assign ram_c_20_0_rdata = ram_c_20_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_c_20_0_enable) begin
      if(ram_c_20_0_wenable) begin
        mem[ram_c_20_0_addr] <= ram_c_20_0_wdata;
        ram_c_20_0_rdata_out <= ram_c_20_0_wdata;
      end else begin
        ram_c_20_0_rdata_out <= mem[ram_c_20_0_addr];
      end
    end 
  end


endmodule



module ram_c_21
(
  input CLK,
  input [20-1:0] ram_c_21_0_addr,
  output [32-1:0] ram_c_21_0_rdata,
  input [32-1:0] ram_c_21_0_wdata,
  input ram_c_21_0_wenable,
  input ram_c_21_0_enable
);

  reg [32-1:0] ram_c_21_0_rdata_out;
  assign ram_c_21_0_rdata = ram_c_21_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_c_21_0_enable) begin
      if(ram_c_21_0_wenable) begin
        mem[ram_c_21_0_addr] <= ram_c_21_0_wdata;
        ram_c_21_0_rdata_out <= ram_c_21_0_wdata;
      end else begin
        ram_c_21_0_rdata_out <= mem[ram_c_21_0_addr];
      end
    end 
  end


endmodule



module ram_c_22
(
  input CLK,
  input [20-1:0] ram_c_22_0_addr,
  output [32-1:0] ram_c_22_0_rdata,
  input [32-1:0] ram_c_22_0_wdata,
  input ram_c_22_0_wenable,
  input ram_c_22_0_enable
);

  reg [32-1:0] ram_c_22_0_rdata_out;
  assign ram_c_22_0_rdata = ram_c_22_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_c_22_0_enable) begin
      if(ram_c_22_0_wenable) begin
        mem[ram_c_22_0_addr] <= ram_c_22_0_wdata;
        ram_c_22_0_rdata_out <= ram_c_22_0_wdata;
      end else begin
        ram_c_22_0_rdata_out <= mem[ram_c_22_0_addr];
      end
    end 
  end


endmodule



module ram_c_23
(
  input CLK,
  input [20-1:0] ram_c_23_0_addr,
  output [32-1:0] ram_c_23_0_rdata,
  input [32-1:0] ram_c_23_0_wdata,
  input ram_c_23_0_wenable,
  input ram_c_23_0_enable
);

  reg [32-1:0] ram_c_23_0_rdata_out;
  assign ram_c_23_0_rdata = ram_c_23_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_c_23_0_enable) begin
      if(ram_c_23_0_wenable) begin
        mem[ram_c_23_0_addr] <= ram_c_23_0_wdata;
        ram_c_23_0_rdata_out <= ram_c_23_0_wdata;
      end else begin
        ram_c_23_0_rdata_out <= mem[ram_c_23_0_addr];
      end
    end 
  end


endmodule



module ram_c_24
(
  input CLK,
  input [20-1:0] ram_c_24_0_addr,
  output [32-1:0] ram_c_24_0_rdata,
  input [32-1:0] ram_c_24_0_wdata,
  input ram_c_24_0_wenable,
  input ram_c_24_0_enable
);

  reg [32-1:0] ram_c_24_0_rdata_out;
  assign ram_c_24_0_rdata = ram_c_24_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_c_24_0_enable) begin
      if(ram_c_24_0_wenable) begin
        mem[ram_c_24_0_addr] <= ram_c_24_0_wdata;
        ram_c_24_0_rdata_out <= ram_c_24_0_wdata;
      end else begin
        ram_c_24_0_rdata_out <= mem[ram_c_24_0_addr];
      end
    end 
  end


endmodule



module ram_c_25
(
  input CLK,
  input [20-1:0] ram_c_25_0_addr,
  output [32-1:0] ram_c_25_0_rdata,
  input [32-1:0] ram_c_25_0_wdata,
  input ram_c_25_0_wenable,
  input ram_c_25_0_enable
);

  reg [32-1:0] ram_c_25_0_rdata_out;
  assign ram_c_25_0_rdata = ram_c_25_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_c_25_0_enable) begin
      if(ram_c_25_0_wenable) begin
        mem[ram_c_25_0_addr] <= ram_c_25_0_wdata;
        ram_c_25_0_rdata_out <= ram_c_25_0_wdata;
      end else begin
        ram_c_25_0_rdata_out <= mem[ram_c_25_0_addr];
      end
    end 
  end


endmodule



module ram_c_26
(
  input CLK,
  input [20-1:0] ram_c_26_0_addr,
  output [32-1:0] ram_c_26_0_rdata,
  input [32-1:0] ram_c_26_0_wdata,
  input ram_c_26_0_wenable,
  input ram_c_26_0_enable
);

  reg [32-1:0] ram_c_26_0_rdata_out;
  assign ram_c_26_0_rdata = ram_c_26_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_c_26_0_enable) begin
      if(ram_c_26_0_wenable) begin
        mem[ram_c_26_0_addr] <= ram_c_26_0_wdata;
        ram_c_26_0_rdata_out <= ram_c_26_0_wdata;
      end else begin
        ram_c_26_0_rdata_out <= mem[ram_c_26_0_addr];
      end
    end 
  end


endmodule



module ram_c_27
(
  input CLK,
  input [20-1:0] ram_c_27_0_addr,
  output [32-1:0] ram_c_27_0_rdata,
  input [32-1:0] ram_c_27_0_wdata,
  input ram_c_27_0_wenable,
  input ram_c_27_0_enable
);

  reg [32-1:0] ram_c_27_0_rdata_out;
  assign ram_c_27_0_rdata = ram_c_27_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_c_27_0_enable) begin
      if(ram_c_27_0_wenable) begin
        mem[ram_c_27_0_addr] <= ram_c_27_0_wdata;
        ram_c_27_0_rdata_out <= ram_c_27_0_wdata;
      end else begin
        ram_c_27_0_rdata_out <= mem[ram_c_27_0_addr];
      end
    end 
  end


endmodule



module ram_c_28
(
  input CLK,
  input [20-1:0] ram_c_28_0_addr,
  output [32-1:0] ram_c_28_0_rdata,
  input [32-1:0] ram_c_28_0_wdata,
  input ram_c_28_0_wenable,
  input ram_c_28_0_enable
);

  reg [32-1:0] ram_c_28_0_rdata_out;
  assign ram_c_28_0_rdata = ram_c_28_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_c_28_0_enable) begin
      if(ram_c_28_0_wenable) begin
        mem[ram_c_28_0_addr] <= ram_c_28_0_wdata;
        ram_c_28_0_rdata_out <= ram_c_28_0_wdata;
      end else begin
        ram_c_28_0_rdata_out <= mem[ram_c_28_0_addr];
      end
    end 
  end


endmodule



module ram_c_29
(
  input CLK,
  input [20-1:0] ram_c_29_0_addr,
  output [32-1:0] ram_c_29_0_rdata,
  input [32-1:0] ram_c_29_0_wdata,
  input ram_c_29_0_wenable,
  input ram_c_29_0_enable
);

  reg [32-1:0] ram_c_29_0_rdata_out;
  assign ram_c_29_0_rdata = ram_c_29_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_c_29_0_enable) begin
      if(ram_c_29_0_wenable) begin
        mem[ram_c_29_0_addr] <= ram_c_29_0_wdata;
        ram_c_29_0_rdata_out <= ram_c_29_0_wdata;
      end else begin
        ram_c_29_0_rdata_out <= mem[ram_c_29_0_addr];
      end
    end 
  end


endmodule



module ram_c_30
(
  input CLK,
  input [20-1:0] ram_c_30_0_addr,
  output [32-1:0] ram_c_30_0_rdata,
  input [32-1:0] ram_c_30_0_wdata,
  input ram_c_30_0_wenable,
  input ram_c_30_0_enable
);

  reg [32-1:0] ram_c_30_0_rdata_out;
  assign ram_c_30_0_rdata = ram_c_30_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_c_30_0_enable) begin
      if(ram_c_30_0_wenable) begin
        mem[ram_c_30_0_addr] <= ram_c_30_0_wdata;
        ram_c_30_0_rdata_out <= ram_c_30_0_wdata;
      end else begin
        ram_c_30_0_rdata_out <= mem[ram_c_30_0_addr];
      end
    end 
  end


endmodule



module ram_c_31
(
  input CLK,
  input [20-1:0] ram_c_31_0_addr,
  output [32-1:0] ram_c_31_0_rdata,
  input [32-1:0] ram_c_31_0_wdata,
  input ram_c_31_0_wenable,
  input ram_c_31_0_enable
);

  reg [32-1:0] ram_c_31_0_rdata_out;
  assign ram_c_31_0_rdata = ram_c_31_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_c_31_0_enable) begin
      if(ram_c_31_0_wenable) begin
        mem[ram_c_31_0_addr] <= ram_c_31_0_wdata;
        ram_c_31_0_rdata_out <= ram_c_31_0_wdata;
      end else begin
        ram_c_31_0_rdata_out <= mem[ram_c_31_0_addr];
      end
    end 
  end


endmodule



module ram_x
(
  input CLK,
  input [20-1:0] ram_x_0_addr,
  output [32-1:0] ram_x_0_rdata,
  input [32-1:0] ram_x_0_wdata,
  input ram_x_0_wenable,
  input ram_x_0_enable
);

  reg [32-1:0] ram_x_0_rdata_out;
  assign ram_x_0_rdata = ram_x_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_x_0_enable) begin
      if(ram_x_0_wenable) begin
        mem[ram_x_0_addr] <= ram_x_0_wdata;
        ram_x_0_rdata_out <= ram_x_0_wdata;
      end else begin
        ram_x_0_rdata_out <= mem[ram_x_0_addr];
      end
    end 
  end


endmodule



module ram_y
(
  input CLK,
  input [20-1:0] ram_y_0_addr,
  output [32-1:0] ram_y_0_rdata,
  input [32-1:0] ram_y_0_wdata,
  input ram_y_0_wenable,
  input ram_y_0_enable
);

  reg [32-1:0] ram_y_0_rdata_out;
  assign ram_y_0_rdata = ram_y_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_y_0_enable) begin
      if(ram_y_0_wenable) begin
        mem[ram_y_0_addr] <= ram_y_0_wdata;
        ram_y_0_rdata_out <= ram_y_0_wdata;
      end else begin
        ram_y_0_rdata_out <= mem[ram_y_0_addr];
      end
    end 
  end


endmodule



module ram_z
(
  input CLK,
  input [20-1:0] ram_z_0_addr,
  output [32-1:0] ram_z_0_rdata,
  input [32-1:0] ram_z_0_wdata,
  input ram_z_0_wenable,
  input ram_z_0_enable
);

  reg [32-1:0] ram_z_0_rdata_out;
  assign ram_z_0_rdata = ram_z_0_rdata_out;
  reg [32-1:0] mem [0:1048576-1];

  always @(posedge CLK) begin
    if(ram_z_0_enable) begin
      if(ram_z_0_wenable) begin
        mem[ram_z_0_addr] <= ram_z_0_wdata;
        ram_z_0_rdata_out <= ram_z_0_wdata;
      end else begin
        ram_z_0_rdata_out <= mem[ram_z_0_addr];
      end
    end 
  end


endmodule

